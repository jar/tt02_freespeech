module jar_pi
(
	input  [7:0] io_in,
	output [7:0] io_out
);
	wire       clk      = io_in[0];
	wire       reset    = io_in[1];
//	wire       stream   = io_in[2];
//	wire [4:0] io_index = io_in[7:3];

	reg [9:0] index;
	//reg [7:0] led_out;
	wire [3:0] code;
	//assign io_out[7:0] = led_out;

	wire j = index[9];
	wire i = index[8];
	wire h = index[7];
	wire g = index[6];
	wire f = index[5];
	wire e = index[4];
	wire d = index[3];
	wire c = index[2];
	wire b = index[1];
	wire a = index[0];

	always @(posedge clk) begin
		if (reset) begin
//			index <= {io_index, index[9:5]};
			index <= 10'b0000000000;
		end
		else begin
//		else if (stream) begin
			index <= index + 1;
//		end

code[3]<=j?(i?(h?((g&!f&e&d&b&a)|(g&f&!d&c&b&a)|(g&!f&e&!d&!b&a)|(g&d&c&!b&a)|(!e&d&!c&!a)|(!f&d&c&!b&a)|(!g&f&!e&d&c)|(f&d&!c&a)|(!f&e&c&!b)|(!g&f&c&!b)|(!g&!d&a)):((g&f&e&!d&!b&!a)|(!g&!f&!d&c&a)|(f&!e&!d&c&b)|(d&!c&b&a)|(!g&!f&!d&!c&!a)|(!g&!e&!c&b&!a)|(!g&!e&d&b&a)|(f&!e&d&!b&!a)|(!d&!c&b&!a)|(g&!e&!b&a)|(!d&!c&!b&a)|(e&d&c&a))):(h?((g&!f&!e&d&b&a)|(!f&!e&d&c&b&a)|(!g&e&!d&!c&b&a)|(!g&e&d&!c&b&!a)|(g&f&!d&!c&b&a)|(!g&f&e&!d&b&!a)|(!g&f&!e&c&b&a)|(!f&!e&!d&!c&b)|(g&f&e&!c&b)|(f&!d&c&!b&a)|(g&f&!e&c&!b)|(g&e&d&c&!b)|(g&f&e&d&c)|(g&!f&e&!a)|(!g&d&!c&!b)|(!g&!e&!d&!a)):((!g&f&d&!c&b&!a)|(!g&!f&e&!d&!c&!a)|(!g&!f&e&d&b&a)|(f&e&c&!b&a)|(!f&!d&c&b&!a)|(g&!f&d&c&a)|(!f&!e&d&!c&b)|(!g&!e&!d&c&b)|(g&f&d&!a)|(g&e&!d&!c)))):(i?(h?((g&e&!d&c&b&!a)|(f&d&!c&b&!a)|(!f&!e&!c&!b&!a)|(!g&f&!e&!d&a)|(!f&!d&c&!b&a)|(f&e&d&!b&a)|(!g&!f&e&d&c)|(g&f&d&!c&!b)|(g&!d&b&a)|(g&d&c&!b)|(g&e&!c&a)|(g&!c&b&!a)|(!g&e&!c&!a)):((g&!f&!e&!c&!b&a)|(g&f&!e&!d&!c&!a)|(f&!e&!d&c&b&a)|(!g&!f&!c&!b&!a)|(!f&!e&c&!b&!a)|(!g&f&e&b&!a)|(g&!f&d&c&a)|(e&!d&c&b&!a)|(!g&e&d&c&!b)|(g&f&!d&!b)|(!f&!d&!c&a)|(!g&e&c&b))):(h?((!f&e&!d&c&!b&!a)|(g&!f&!e&!c&!b&!a)|(g&f&e&d&!c&!a)|(!f&e&c&b&a)|(!g&!d&c&b&a)|(!f&e&!c&!b&a)|(!f&!e&b&!a)|(f&d&c&!b)|(!g&f&e&c)|(!e&!c&b&!a)|(g&!e&!b&a)):((!g&!f&!e&c&b&!a)|(g&f&!e&!d&!b&a)|(g&e&!d&!c&!a)|(g&!e&!d&c&!a)|(f&!e&d&b&!a)|(!f&!e&d&b&a)|(!g&f&!e&b&a)|(!g&!f&e&b&a)|(g&!f&e&!b&a)|(!g&!f&!e&!b&a)|(!g&f&!c&!b&!a)|(f&e&d&a)|(!g&f&c&!b)|(d&c&!b&!a))));

code[2]<=j?(i?(h?((!g&!f&!e&!d&!c&!b&a)|(g&f&!e&d&c&b&!a)|(!g&!f&e&d&!c&!b&!a)|(g&f&e&d&!b&!a)|(g&f&!e&!d&!c&b)|(!g&!f&d&c&b&a)|(!g&f&!e&d&c&!b)|(!f&e&!d&c&!b&a)|(g&!f&!e&d&!c&b)|(!g&f&e&d&!c&b&a)|(!g&f&e&!d&c&b&!a)|(!g&!e&!d&!c&b&!a)|(!g&f&e&!d&c&!b&a)|(!g&!f&e&!d&b&!a)|(!g&!e&d&!c&b&!a)|(f&e&d&!c&b&!a)|(!g&f&!e&d&!c&!a)|(!f&e&d&c&!b&!a)|(!g&!f&e&d&c&!a)|(f&e&d&c&b&a)|(!g&!f&!e&!d&b&!a)|(g&e&!d&c&b)|(!g&d&c&!b&!a)|(!g&!f&e&!d&!c&b)|(g&!f&!d&b&a)|(!g&e&c&!b&!a)|(f&e&!d&!c&!b)):((!g&!f&!e&d&c&b&a)|(!g&f&e&d&c&b&a)|(!g&f&!e&d&c&b&!a)|(!g&!f&e&!d&!c&!b&a)|(!g&f&!e&!d&c&b&a)|(!g&!f&!e&d&c&!b&!a)|(!g&f&e&d&!c&!b&!a)|(!g&f&!d&c&b&!a)|(g&!f&!e&d&!c&a)|(g&f&e&c&!b&!a)|(!g&f&!e&!d&!c&!a)|(g&f&e&d&!c&a)|(g&f&!e&d&!c&!a)|(!g&f&!d&c&!b&a)|(!g&!f&d&!c&!b&a)|(!g&f&!e&d&!b&a)|(!g&!f&!e&!d&!c&b&a)|(g&!f&!d&c&!b&!a)|(g&f&!d&c&b&a)|(g&e&d&c&b&!a)|(!g&!f&e&c&!b&!a)|(g&f&e&d&c&!b)|(!f&!e&!d&c&b&!a)|(g&!e&!d&!c&b)|(f&!e&d&!c&b))):(h?((g&f&e&d&!c&b&!a)|(!g&!f&!e&d&c&!b&a)|(!g&f&!e&!c&!b&a)|(g&f&!e&d&!c&!b&!a)|(g&!f&e&!d&!c&!b&!a)|(!g&f&e&!d&!c&b&!a)|(g&!f&e&!d&b&a)|(!g&f&e&d&c&!b&a)|(!g&f&e&d&!c&!b&!a)|(!g&f&e&!d&c&!b&!a)|(g&f&e&!d&!c&!b&!a)|(!g&!f&e&!d&!c&!b)|(g&!f&!d&c&!b&!a)|(!g&f&d&c&b&!a)|(!g&!f&!e&!d&c&!a)|(g&f&!e&c&b&!a)|(g&e&!d&!c&b&a)|(g&f&!d&c&!b&a)|(f&!e&!d&!c&!b&a)|(!f&e&d&!b&!a)|(!g&!f&d&!c&!a)|(!g&f&!e&d&c&!a)|(g&!e&!d&c&!b)|(!g&f&!e&!d&!c)|(!g&!f&!e&b&!a)|(f&!e&!d&c&a)):((!g&!f&e&!d&c&!b&!a)|(!g&!f&!e&!d&c&b&!a)|(g&f&!e&!d&c&!b)|(!g&f&d&!c&!b&!a)|(g&e&d&c&b&!a)|(g&f&!e&c&b&a)|(g&!e&d&c&b&a)|(g&!e&d&!c&!b&a)|(!f&e&d&c&!b&a)|(g&e&!d&b&!a)|(g&!e&d&b&!a)|(g&!f&e&!d&!a)|(g&f&e&d&!c)|(!g&d&!c&b&a)|(!f&!e&!d&b&a)|(!g&e&d&!c&b)|(!f&!d&!c&!b&a)|(!g&!f&!d&b&a)|(g&!f&!e&!c&!b)|(!g&!f&!e&!d&!b)|(!g&f&e&!c&!b&!a)|(!g&f&!d&!c&!b&a)|(!g&f&!e&c&!b&a)|(f&e&!d&!c&a)|(g&!d&!c&b&!a)))):(i?(h?((g&e&d&!c&b&a)|(g&!f&!e&d&!c&!b&!a)|(!g&f&!e&d&!c&b&a)|(!g&!f&!e&!d&c&!b&!a)|(g&!e&!d&c&b&a)|(g&!f&!e&!d&b&!a)|(g&!e&!d&!c&!b&a)|(g&f&e&d&b&!a)|(g&f&e&!c&b&!a)|(!g&e&d&!c&!b&!a)|(!g&!e&d&c&b&!a)|(!g&f&!e&!d&!b&!a)|(g&!f&!e&!d&!b&a)|(g&!f&e&!d&!b&!a)|(!g&!f&e&c&b&!a)|(!f&!e&c&b&!a)|(!g&!f&!e&!c&a)|(!f&d&!c&b&a)|(!g&e&c&!b&a)|(!f&e&!d&!b&a)|(!f&e&d&c&!b)|(g&!f&e&b&a)):((!g&!f&!e&d&!c&!b&!a)|(g&!f&!e&!d&!c&!b&a)|(!g&!f&e&!d&c&!b&a)|(g&!f&!e&!d&c&b&!a)|(!g&f&e&d&c&!b)|(g&f&e&d&!c&a)|(!g&f&!e&c&b&!a)|(g&!f&e&d&c&a)|(!f&!e&!d&!c&b&!a)|(!g&!f&e&!d&b&!a)|(!g&!f&!e&!c&b&a)|(g&e&d&!c&b&!a)|(!g&!f&!d&c&b&a)|(g&!f&e&d&!c&!b&!a)|(!g&f&e&!d&!c&b&a)|(g&f&!e&!d&!b&!a)|(g&f&!d&!c&!b&!a)|(g&f&!e&!c&!b&!a)|(!g&f&!e&d&c&!a)|(!f&!e&d&c&!b&a)|(!g&f&!e&!d&!c&a)|(!g&f&e&!d&c&b)|(!f&e&d&c&b&a)|(g&e&!d&!c&b&a)|(!g&f&!c&!b&a)|(!g&e&!d&!c&!b)|(g&e&c&!b&!a)|(!g&!d&!c&!b&a))):(h?((!g&!f&!e&!d&!c&!b&!a)|(!g&f&e&d&!c&!b&a)|(g&f&e&!d&!c&!b&!a)|(g&f&!e&!d&!c&b&!a)|(!g&!f&e&d&c&b)|(!g&f&d&c&!b&a)|(g&f&!e&c&!b&!a)|(!g&!f&e&!d&!c&!a)|(!g&f&e&!d&c&!a)|(!g&e&d&!c&!b&!a)|(g&!f&e&!d&c&!b)|(!g&!e&!d&!c&b&a)|(!g&!f&e&d&c&!b&a)|(g&!f&e&c&!b&!a)|(g&!f&e&!d&b&!a)|(g&f&!d&!c&b&a)|(!g&f&e&!d&!c&b)|(g&f&!d&!c&!b&a)|(!g&f&!d&b&a)|(g&!f&d&!c&b)|(g&e&!d&!c&b&a)|(g&f&e&d&c)|(g&!e&d&!c&a)|(g&!e&!d&!c&!b)|(!g&!f&!e&c&!a)):((g&!f&e&d&c&!b&a)|(g&!f&!e&!d&c&b&!a)|(g&!f&!e&d&c&!b&!a)|(g&!f&!e&!d&b&a)|(g&!f&e&!c&b&a)|(g&f&d&c&b&!a)|(!g&f&!d&!c&!b&!a)|(!g&f&d&!c&b&!a)|(!g&!f&e&!d&c&a)|(g&f&e&d&!c&!b)|(!g&!f&!e&!c&b&a)|(g&f&!e&!d&c&!b&!a)|(!g&!e&!d&c&!b&a)|(!g&e&!d&c&!b&!a)|(!g&e&d&c&b&!a)|(!f&!e&d&!c&!b&a)|(g&f&!e&d&!b&a)|(!f&e&d&!c&!b&!a)|(!g&f&e&d&c&!b)|(g&f&!e&!d&!c&a)|(!g&!f&d&c&b&!a)|(!g&f&e&!c&!b&a)|(!g&!e&d&!c&!b&!a)|(g&f&e&c&b))));

code[1]<=j?(i?(h?((g&f&e&!d&!c&!b&a)|(g&!f&!d&c&a)|(!g&!f&e&d&c&b&a)|(!g&!f&e&d&!c&!b&!a)|(g&!f&!e&c&!b&a)|(g&f&!e&!d&!b&!a)|(!g&f&!e&d&!c&!b&a)|(g&!f&!e&!d&!c&!b)|(f&!e&d&c&b&a)|(!g&!f&!e&!d&c&!b&a)|(!g&f&d&c&!b&!a)|(!g&!f&d&!c&!b&a)|(!g&e&!d&!c&!b&!a)|(g&!f&!e&d&!c&b)|(!g&f&e&d&!c&b&a)|(!g&f&e&!d&c&b&!a)|(!g&!e&!d&!c&b&!a)|(!g&f&e&!d&c&!b&a)|(!g&!f&e&!d&b&!a)|(f&!e&d&!c&b&!a)|(g&e&!d&b&!a)|(g&f&e&d&c)|(!g&!f&!e&!c&b&a)|(g&!f&!d&c&b)|(f&!e&!d&!c&!a)|(!g&f&!e&!d&b)|(g&!f&!d&b&a)):((!g&f&!e&d&c&b&!a)|(g&!f&!e&!c&!b&!a)|(g&!f&d&!c&b&a)|(!g&f&e&d&b&!a)|(!g&!f&!e&!d&!c&b&a)|(g&!f&!d&c&!b&!a)|(g&f&!d&c&b&a)|(g&e&d&c&b&!a)|(!g&!f&e&c&!b&!a)|(g&!f&!e&!d&!c&!b)|(g&f&e&d&c&!b)|(!g&e&!d&!c&b&!a)|(g&f&!e&!d&!c&!a)|(g&f&e&!c&!b&a)|(!f&e&d&c&!b&a)|(g&f&!e&d&c&!b)|(!g&!f&!d&b&!a)|(g&!e&d&b&!a)|(!g&!f&e&!b&a)|(f&e&!d&c&a)|(!g&!d&c&!b&!a)|(f&!e&c&!b&!a)|(f&e&d&!c&a))):(h?((!g&!f&e&d&c&!b&a)|(g&f&e&d&!c&!b&a)|(g&!f&e&!d&!c&!b&!a)|(!g&f&e&!d&!c&b&!a)|(!g&e&d&!c&b&a)|(!g&f&e&d&c&!b&!a)|(!g&f&e&!d&c&!b&!a)|(!g&!f&e&!d&c&b)|(g&e&!d&c&b&!a)|(g&!f&!e&c&!b&a)|(!g&f&e&c&b&a)|(f&!e&d&c&b&!a)|(g&f&!e&!d&c&a)|(!g&f&e&!d&!c&!b)|(!g&!f&!e&!d&c&!b)|(g&e&!d&!c&b&a)|(g&f&!d&c&!b&a)|(f&!e&!d&!c&!b&a)|(!g&f&!e&d&!c&!b)|(!f&!e&d&!c&!a)|(!g&!f&!e&!c&b)|(g&f&!e&!d&!b&!a)|(g&f&!e&!c&!a)|(!g&!f&!e&b&!a)):((!g&!f&e&!d&c&!b&!a)|(!g&!f&!e&!d&c&b&!a)|(!g&!f&!e&d&!c&!b&!a)|(g&f&e&!d&c&a)|(f&!e&!d&!c&!b&a)|(!g&e&d&!c&b&a)|(!g&!f&!e&d&b&a)|(!g&!e&!d&!c&b&a)|(!g&f&d&!c&!b&!a)|(g&e&d&c&b&!a)|(g&f&!e&c&b&a)|(!g&f&e&d&b&!a)|(g&f&d&!c&!b&!a)|(g&!e&d&c&b&a)|(!g&f&!e&d&c&!b)|(!g&!f&e&d&c&!b)|(g&f&!e&b&!a)|(!g&f&e&c&!a)|(f&!e&d&c&a)|(!f&e&d&!c&!b)|(!g&!f&c&!b&a)|(g&!f&!e&!d&!b)|(!g&f&e&!c&!b&!a)|(!g&f&!d&!c&!b&a)|(!g&f&!e&c&!b&a)|(g&!d&!c&b&!a)|(g&f&e&!c&b)|(g&!f&!c&!b)))):(i?(h?((f&!d&c&!b&a)|(g&f&!e&!d&!c&!b&!a)|(!g&!f&e&d&c&!b&a)|(!g&f&!e&d&!c&b&a)|(!g&!f&!e&!d&c&!b&!a)|(g&f&!e&!d&c&b)|(!g&f&e&!d&c&!b)|(!g&f&d&!c&!b&!a)|(!g&!e&d&c&b&!a)|(!g&f&!e&d&c&b)|(!g&e&!d&!c&b&a)|(g&!f&e&!d&!b&!a)|(g&!d&c&!b&a)|(g&!f&d&c&b)|(g&!f&!e&d&!c)|(!g&!f&e&!d&b)|(g&!f&e&c&!a)|(!g&!f&e&!c&b)|(g&f&d&!b&a)|(!g&e&d&!c&!a)|(g&f&e&d)):((!g&!f&!e&d&!c&!b&!a)|(g&f&e&!d&!c&!b&a)|(g&!f&!e&!d&!c&!b&a)|(!g&!f&e&!d&c&!b&a)|(g&f&d&c&!b&a)|(!g&f&!e&d&b&a)|(!g&e&d&!c&!b&a)|(!f&!e&d&!c&b&!a)|(f&e&d&!c&b&!a)|(g&!f&e&!d&!c&!a)|(f&!e&!d&!c&b&a)|(g&!e&d&c&b&!a)|(!g&!f&!d&c&b&!a)|(f&e&!d&c&b&a)|(g&!e&!d&c&b&a)|(g&!f&e&d&!c&!b&!a)|(!g&f&e&!d&!c&b&a)|(g&f&!e&!c&!b&!a)|(!g&f&!e&d&c&!a)|(!f&!e&d&c&!b&a)|(!g&f&!e&!d&!c&a)|(!g&f&e&!d&c&b)|(!g&!f&e&!c&b&a)|(!f&e&d&c&b&a)|(!g&!e&c&!b&a)|(!f&e&d&c&!a)|(!g&!f&e&c&!a)|(!g&!e&!d&!c&b)|(g&e&d&b&a))):(h?((!g&!f&!e&!d&!c&!b&!a)|(!g&f&e&d&!c&!b&a)|(g&f&e&!d&!c&!b&!a)|(g&!f&!e&!d&c&!b&a)|(!g&!f&!e&d&!c&!a)|(!g&!f&!e&d&c&a)|(!f&!e&d&c&!b&!a)|(!f&!e&d&!c&!b&a)|(f&!e&d&!c&b&a)|(!g&f&e&d&!c&b)|(g&e&d&c&b&!a)|(!g&e&!d&c&b&!a)|(f&!e&!d&!c&!b&a)|(g&e&!d&!c&b&!a)|(g&!e&!d&!c&b&a)|(g&e&!d&c&!b&a)|(!g&!f&e&d&c&!b&a)|(g&f&!e&d&c&!a)|(g&!f&e&c&!b&!a)|(g&f&!d&!c&b&a)|(g&f&!e&d&!c&!b)|(f&!e&!d&c&b&a)|(g&!f&e&d&!c&!b)|(f&!e&c&b&!a)):((!g&f&!e&d&c&b&a)|(g&!f&!e&!d&c&b&!a)|(g&!f&!e&d&c&!b&!a)|(g&f&e&!d&!c&!b)|(f&e&!d&c&b&!a)|(!g&!f&!d&c&b&a)|(!g&f&!e&!c&b&!a)|(g&f&!e&!d&c&!b&!a)|(!g&e&!d&!c&!b&!a)|(g&!e&d&c&!b&a)|(f&e&d&!c&!b&a)|(g&!f&!e&d&!b&a)|(g&f&!e&!d&!c&a)|(g&!f&!e&!d&!c&a)|(!g&!f&d&c&b&!a)|(!g&!e&d&!c&!b&!a)|(!f&e&d&c&!b&!a)|(!g&f&!e&d&!b&!a)|(g&f&!d&b&a)|(g&e&!d&b&a)|(!f&!e&!d&!c&!b)|(!f&d&!c&b&!a)|(g&e&c&!b&!a)|(!f&e&d&b&!a)|(!g&!f&e&b&!a)|(!g&!f&e&!b&a))));

code[0]<=j?(i?(h?((g&f&!e&d&c&b&!a)|(!g&f&!e&d&!c&!b&a)|(g&!f&!e&c&!b&!a)|(!g&!f&!e&!d&c&!b&a)|(g&f&!e&!c&!b&a)|(g&f&!e&!d&c&b)|(g&!f&e&d&b&a)|(g&f&!d&c&b&a)|(g&!f&e&!d&!b&a)|(!g&f&e&d&!c&b&a)|(!g&f&e&!d&c&b&!a)|(!g&f&e&!d&c&!b&a)|(f&!e&d&!c&b&!a)|(!g&!e&d&!c&b&!a)|(f&e&d&!c&b&!a)|(!g&f&!e&d&!c&!a)|(!f&e&d&c&!b&!a)|(!g&!f&e&d&c&!a)|(f&e&d&c&b&a)|(!g&!f&!e&!c&b&a)|(!g&!f&!e&!d&b&!a)|(!g&!f&e&!d&!c&b)|(g&!f&e&!c&!b)|(!f&!e&!d&!c&!a)|(!g&f&e&!c&!a)|(f&e&!d&!b&!a)|(!f&!d&!c&b&a)|(!g&!e&!d&b&a)|(!g&!d&!c&b&a)|(g&d&c&!b&a)|(!f&d&c&!b&a)|(!g&f&!e&d&c)|(!g&e&c&!b&!a)|(f&e&!d&!c&!b)|(!f&e&d&!c)):((!g&!f&e&!d&!c&!b&a)|(!g&f&!e&!d&c&b&a)|(!g&!f&!e&d&c&!b&!a)|(!g&f&e&d&!c&!b&!a)|(g&!f&e&!d&c&a)|(!g&!f&e&!c&!b&!a)|(!f&e&d&c&b&!a)|(!g&f&!e&!d&!c&!b)|(!g&!f&!e&!d&!c&b&a)|(g&!f&!e&!d&!c&!b)|(!g&e&!d&!c&b&!a)|(!f&!e&!d&c&b&!a)|(g&f&!e&!d&!c&!a)|(g&f&e&!c&!b&a)|(!f&e&d&c&!b&a)|(g&f&!e&d&c&!b)|(!f&e&!c&b&a)|(!f&e&!d&!b&!a)|(g&!f&!e&d&c)|(g&f&!c&b&a)|(g&!f&!e&d&!b)|(g&f&e&d&!c)|(!g&!f&c&!b&a)|(f&e&d&b&a)|(g&d&c&!b&!a)|(!g&!f&!d&!c&!a)|(!g&!e&!c&b&!a)|(!g&!e&d&b&a)|(f&!e&d&!b&!a)|(f&!e&d&!c&b))):(h?((!g&f&e&d&c&!b&a)|(!g&f&e&d&!c&!b&!a)|(!g&f&e&d&c&!b&!a)|(g&f&e&!d&!c&!b&!a)|(g&!f&!d&c&b&!a)|(!g&!f&!d&c&!b&a)|(!g&e&!d&!c&b&a)|(g&!e&!d&c&!b&!a)|(!g&e&d&!c&b&!a)|(g&f&!d&!c&b&a)|(!g&f&e&!d&b&!a)|(!g&f&!e&c&b&a)|(!g&f&!e&d&!c&!b)|(g&!f&!e&!c&a)|(g&f&!e&!d&!b&!a)|(!g&f&!e&d&c&!a)|(g&!f&!e&c&b)|(!g&!e&!c&b&!a)|(!g&!f&!e&!d&!c)|(!g&!e&d&!b&!a)|(f&!e&d&!c&!a)|(g&e&d&c&!b)|(f&!e&c&!b&!a)|(g&f&e&d&c)|(!f&e&d&a)|(f&!e&!d&c&a)|(g&f&e&a)|(!f&!e&!d&b)|(g&f&d&!b)):((g&!f&!e&d&c&!b&!a)|(!g&!e&!d&c&!b&!a)|(!g&!f&!e&d&!c&!b&!a)|(g&!f&e&!c&!b&!a)|(!g&f&!e&!d&c&!a)|(g&f&!e&d&c&b)|(g&!e&!d&c&!b&a)|(!g&f&d&!c&b&!a)|(!g&!f&e&!d&!c&!a)|(!g&!f&e&d&b&a)|(!g&f&e&d&b&!a)|(g&f&d&!c&!b&!a)|(g&!e&d&!c&!b&a)|(!f&e&d&c&!b&a)|(!g&f&!e&d&c&!b)|(!g&!f&e&d&c&!b)|(g&!e&!d&!c&!a)|(g&!d&!c&b&a)|(f&e&!d&c&!b)|(!f&e&!d&c&b)|(!g&!f&d&c&b)|(!g&f&e&!c&!b&!a)|(!g&f&!d&!c&!b&a)|(!g&f&!e&c&!b&a)|(f&e&!d&!c&a)|(g&f&e&!c&b)|(f&e&!b&a)|(!g&e&c&a)))):(i?(h?((!g&!f&!e&!d&c&b)|(g&f&!d&c&!b&!a)|(!g&!f&d&!b&!a)|(!g&f&!e&d&c&b)|(g&e&!d&c&b&!a)|(!g&f&!e&!d&!b&!a)|(g&!f&!e&!d&!b&a)|(!g&e&!d&!c&b&a)|(!g&!f&e&c&b&!a)|(g&f&!e&b&a)|(!g&f&!e&c&!b)|(!f&!e&d&!c&b)|(!g&!d&!c&b&!a)|(!g&f&!c&!b&a)|(!f&e&!d&!c&!a)|(!g&f&!e&!d&a)|(g&e&d&!b&!a)|(!f&!d&c&!b&a)|(g&e&!c&!b&!a)|(f&e&d&!b&a)|(!g&!f&e&d&c)|(g&f&d&!c&!b)|(g&f&d&!b&a)|(g&!f&e&b&a)|(!g&e&d&!c&!a)|(f&e&!c&a)|(!f&d&c&!b)|(!g&f&e&b)):((g&f&!e&d&!c&b&a)|(g&f&e&d&c&b)|(g&f&e&!d&!c&!b&a)|(g&!f&!e&!d&c&b&!a)|(f&!e&d&c&!b)|(g&!e&d&c&!b&!a)|(g&!e&!d&!c&!b&!a)|(g&!e&!d&c&!b&a)|(!g&!f&!e&!d&c&!a)|(g&!f&e&!d&c&b)|(g&!f&!e&!c&!b&a)|(g&f&!e&!d&!c&!a)|(g&!f&e&d&!c&!b&!a)|(f&!e&!d&c&b&a)|(!g&f&e&!d&!c&b&a)|(g&f&!e&!d&!b&!a)|(g&f&!d&!c&!b&!a)|(!g&!f&e&!c&b&a)|(g&e&!d&!c&b&a)|(!g&f&!e&d&!a)|(g&f&d&c&!a)|(!g&!f&d&b&!a)|(!f&e&d&b&!a)|(g&!f&e&!c&a)|(!g&e&d&!c&b)|(!g&e&d&c&!b)|(!g&!d&!c&!b&a))):(h?((g&f&!e&!d&!c&b&!a)|(g&!f&!e&!d&c&!b&a)|(!g&!e&d&!c&b)|(!g&e&d&c&!b&!a)|(!g&!e&!d&c&!b&!a)|(f&e&!d&c&!b&!a)|(g&f&e&!c&b&a)|(g&e&d&c&!b&a)|(!g&e&!d&!c&!b&!a)|(!f&e&!d&!c&!b&a)|(!g&!f&e&d&c&!b&a)|(!g&e&!d&c&!b&a)|(g&!f&!e&!c&!b&!a)|(g&f&e&d&!c&!a)|(g&f&!e&d&c&!a)|(g&!f&e&!d&b&!a)|(g&f&!e&d&!c&!b)|(f&!e&!d&c&b&a)|(g&!f&e&d&!c&!b)|(!g&f&e&!d&!c&b)|(g&f&!d&!c&!b&a)|(!g&f&!e&d&a)|(g&e&!d&!c&b&a)|(!g&!f&d&!c&b)|(!g&d&c&b&a)|(!f&!e&!d&!c&b)|(g&!e&c&b&a)|(g&!d&c&b&a)|(!g&!f&!e&c&!a)):((g&!f&e&!d&!c&!b)|(g&!f&e&c&b&a)|(g&!f&e&d&b&a)|(!f&!e&!d&c&!b&a)|(g&f&!e&!d&c&!b&!a)|(g&f&e&c&!b&!a)|(g&f&!e&!d&!b&a)|(g&!f&!e&!d&!c&a)|(!g&f&e&!c&!b&a)|(!f&e&d&c&!b&!a)|(!g&f&!e&d&!b&!a)|(!g&e&!d&!c&!a)|(f&!e&d&c&b)|(!g&!f&!c&b&!a)|(!g&!f&!e&!d&!a)|(f&e&d&!c&a)|(!g&f&!e&c&b)|(f&!e&!c&!b&!a)|(f&e&!d&!b&!a)|(!g&d&!c&!b&a)|(!g&f&!c&!b&!a)|(!g&d&c&b)|(!g&!e&d&a))));
		end

	end

	decoder decoder(.code(code), .segments(io_out));

endmodule

module jar_pi
(
	input  [7:0] io_in,
	output [7:0] io_out
);
	wire       clk      = io_in[0];
	//wire       reset    = io_in[1];
	//wire       stream   = io_in[2];
	//wire [4:0] io_index = io_in[7:3];

	reg [9:0] index;
	//reg [7:0] led_out;
	wire [3:0] hex;
	//assign io_out[7:0] = led_out;

	wire v0 = index[9];
	wire v1 = index[8];
	wire v2 = index[7];
	wire v3 = index[6];
	wire v4 = index[5];
	wire v5 = index[4];
	wire v6 = index[3];
	wire v7 = index[2];
	wire v8 = index[1];
	wire v9 = index[0];

	wire n0 = !v0;
	wire n1 = !v1;
	wire n2 = !v2;
	wire n3 = !v3;
	wire n4 = !v4;
	wire n5 = !v5;
	wire n6 = !v6;
	wire n7 = !v7;
	wire n8 = !v8;
	wire n9 = !v9;

	always @(posedge clk) begin
	//	if (reset) begin
	//		index <= {io_index, index[9:5]};
	//	end
	//	else if (stream) begin
			index <= index + 1;
	//	end

hex[3] <= v0 ? ((!v1&!v1&v3&!v4&v5&!v6&!v7&v8&v9) | (!v1&!v1&v3&!v4&!v5&!v6&v7&v8
    &!v9) | (v1&v1&v3&!v4&v5&!v6&v7&!v8&!v9) | (v1&!v1&v3&v4&!v5&!v6&v7
    &v8&!v9) | (!v1&v1&!v3&v4&v5&v6&!v7&v8&!v9) | (v1&v1&!v3&v4&!v5&v6&v7
    &v8&!v9) | (v1&!v1&v3&v4&v5&v6&v7&v8&v9) | (!v1&v1&!v3&!v4&!v5&!v6&!v7
    &!v8&!v9) | (v1&!v1&!v3&!v4&!v5&!v6&v7&!v8&v9) | (v1&v1&v3&v4&!v5&!v6
    &v7&v8&v9) | (!v1&v1&v3&!v4&v5&v6&v8&!v9) | (!v1&!v1&!v3&v4&!v5&v6&!v7
    &v8&!v9) | (v1&v1&v3&!v4&v5&v6&v8&v9) | (v1&!v1&!v3&v4&!v5&v6&v7&v8
    &v9) | (!v1&v1&!v3&v4&!v5&v6&v7&v8&v9) | (v1&!v1&v3&v5&!v6&!v7&v8&!v9) | (
    !v1&v1&v3&v5&!v6&!v7&v8&!v9) | (v1&v3&!v4&v5&!v6&!v7&!v8&v9) | (!v1
    &v3&!v4&!v5&v6&!v7&v8&v9) | (v1&!v1&!v3&v4&!v5&v6&!v7&!v8&!v9) | (v1
    &v3&!v4&v5&v6&v7&!v8&v9) | (!v1&v1&v3&!v4&!v5&!v6&!v7&v8) | (!v1&v1
    &!v4&!v5&v6&v7&v8&v9) | (!v1&v1&v3&v4&v5&v6&v8&v9) | (!v1&v3&!v4&!v5
    &v6&v7&!v8&v9) | (v1&v1&!v4&v5&!v6&!v7&!v8&v9) | (!v1&!v3&!v4&!v5&v6
    &!v7&v8&!v9) | (!v1&v3&v4&v5&!v6&!v7&!v8&!v9) | (v1&v1&!v4&!v5&v6&!v7
    &!v8&!v9) | (v1&!v1&v3&!v5&!v6&v7&!v8&v9) | (!v1&v1&!v3&!v4&v6&!v7&!v8
    &v9) | (!v1&!v1&v4&v5&v6&v7&!v8&v9) | (!v1&v1&!v3&v4&!v6&v7&v8&!v9) | (
    !v1&!v3&v4&v5&!v6&v7&!v8&v9) | (v1&v1&!v3&v4&v5&!v6&v8&v9) | (v1&!v1
    &!v3&!v4&!v5&!v6&!v7&!v8) | (v1&!v1&v3&v4&!v5&!v7&!v8&v9) | (v1&!v3
    &v4&v5&v6&v7&!v8&v9) | (!v1&!v1&!v3&v4&!v5&!v6&v7&v8) | (v1&v1&v4&!v5
    &v6&!v7&v8&v9) | (v1&v1&v3&v4&!v5&v6&!v7&!v8) | (v1&!v1&!v3&v4&!v6&!v7
    &!v8&v9) | (v1&!v3&v4&v5&v6&!v7&!v8&v9) | (v1&!v3&v4&!v5&!v6&v7&!v8
    &!v9) | (v1&v1&!v3&v4&!v5&!v6&!v8&v9) | (!v1&!v1&!v3&!v4&v5&!v6&v8&!v9) | (
    !v1&!v3&!v4&v5&!v6&!v7&!v8&!v9) | (v1&!v1&!v3&!v4&v6&!v7&v8&v9) | (
    !v1&v1&v3&!v5&!v6&!v7&v8&v9) | (!v1&v1&!v3&v5&!v6&!v7&v8&v9) | (v1&v1
    &!v3&!v4&v6&v7&!v8&v9) | (v1&v3&v4&!v5&v6&v7&!v8&v9) | (!v1&!v4&v5&v6
    &v7&v8&v9) | (v1&!v3&!v4&!v6&v7&v8&v9) | (!v1&v3&v4&v6&v7&!v8&!v9) | (
    v1&v1&v3&v4&v6&!v7&v9) | (!v1&v1&v3&v4&v5&v6&v7)) :
    ((v1&!v2&!v3&!v4&v5&v6&!v7&!v8&!v9) | (!v1&!v2&!v3&v4&!v5&v6&v7&v8
    &!v9) | (v1&v2&!v3&v4&v5&v6&!v7&!v8&v9) | (!v1&!v2&!v3&!v4&!v5&!v6&v7
    &v8&!v9) | (!v1&!v2&v3&v4&!v5&!v6&v7&v8&!v9) | (v1&v2&v3&!v4&v5&v6&!v7
    &!v8&v9) | (v1&v2&!v3&!v4&!v5&!v6&v7&!v8&v9) | (v1&!v2&!v3&!v4&v5&v6
    &v7&!v8&v9) | (!v1&!v2&!v3&v4&!v5&!v6&v7&!v8&!v9) | (!v1&v2&!v3&!v4
    &v5&!v6&v7&!v8&!v9) | (!v1&!v2&v3&v4&!v5&v6&v7&!v8&!v9) | (!v1&!v2&!v3
    &!v4&!v5&!v6&!v7&!v8&v9) | (!v1&!v2&v3&v4&v5&v6&v7&!v8&v9) | (v1&!v2
    &v3&v4&!v5&!v6&!v7&v8&!v9) | (v1&v2&!v3&!v4&v5&v6&v7&v8&v9) | (v1&v2
    &!v3&!v4&!v5&v6&!v7&!v8&!v9) | (!v1&!v2&!v3&v4&v5&v6&!v7&!v8&!v9) | (
    v1&!v2&v3&!v4&!v5&v6&!v7&!v8&v9) | (!v1&v2&v3&!v4&!v5&v6&!v7&!v8&!v9) | (
    v1&!v3&v4&v5&!v6&!v7&v8&!v9) | (v1&v2&v3&!v4&v5&!v7&v8&!v9) | (v1&v2
    &v3&v4&!v5&!v6&!v7&v8) | (v1&!v2&!v3&v4&v5&v6&v7&v8) | (v1&v2&!v4&!v5
    &!v6&!v7&!v8&!v9) | (!v1&v3&v4&!v5&v6&!v7&v8&!v9) | (v1&v3&!v4&!v5&!v6
    &!v7&v8&v9) | (v1&v2&v3&v4&v5&!v6&!v7&v9) | (v1&v2&v3&v4&v5&!v6&v7&v8) | (
    v1&v2&v3&v4&!v5&v6&!v8&!v9) | (!v1&!v2&!v3&!v4&v5&!v7&v8&v9) | (!v1
    &v2&v3&!v4&!v5&v7&v8&!v9) | (!v1&v2&!v3&v4&v5&v6&v7&v8) | (v1&!v2&!v3
    &!v4&!v5&!v6&!v8&!v9) | (!v1&!v2&!v3&v4&!v5&!v6&v8&v9) | (!v1&v2&!v3
    &!v5&!v6&!v7&v8&!v9) | (v1&!v2&v3&v5&!v6&v7&v8&!v9) | (!v2&v3&!v4&!v5
    &v6&v7&v8&v9) | (!v1&v2&v3&!v4&v5&v7&v8&v9) | (v1&v2&!v3&v5&!v6&!v7
    &!v8&!v9) | (v1&!v2&v3&v4&!v5&!v6&!v8&v9) | (!v1&v2&!v3&!v4&!v6&v7&v8
    &v9) | (!v1&!v2&v3&!v4&!v5&v6&v8&v9) | (!v2&!v3&!v4&!v5&v6&v7&!v8&!v9) | (
    !v1&v2&!v3&v4&v6&v7&!v8&!v9) | (!v1&v2&!v3&!v4&v5&!v7&!v8&v9) | (!v1
    &!v2&v3&v5&!v6&!v7&v8&!v9) | (v1&!v2&v3&v4&!v6&v7&!v8&v9) | (!v2&v3
    &!v4&!v5&!v6&v7&!v8&!v9) | (!v2&v3&!v4&v5&!v6&!v7&!v8&v9) | (!v1&!v2
    &v3&!v4&v5&!v7&!v8&v9) | (!v1&!v3&v4&v5&!v6&v7&!v8&v9) | (!v1&v3&v4
    &!v5&!v6&v7&!v8&v9) | (!v1&!v2&v3&!v4&v5&!v6&!v8&v9) | (!v1&v2&v3&!v5
    &v6&v7&!v8&v9) | (v1&v2&!v3&v4&!v5&!v6&!v7&v9) | (!v1&v2&!v4&!v5&!v6
    &!v7&v8&!v9) | (v1&!v3&v4&!v5&!v6&v7&v8&v9) | (!v1&!v2&v4&v5&v6&!v7
    &v8&v9) | (!v1&v2&v3&v4&v5&v6&!v7&!v9) | (!v1&!v2&!v3&v4&v6&!v7&v8&v9) | (
    !v1&!v3&v4&v5&v6&v7&v8&v9) | (v1&v3&!v4&!v5&v6&v7&!v8&!v9) | (!v1&!v2
    &!v3&!v4&v6&v7&v8&v9) | (v1&v2&v3&!v4&!v5&v6&v7&!v8) | (!v1&v2&!v4&v5
    &!v6&!v7&!v8&v9) | (!v1&!v2&v3&!v4&v5&!v6&!v7&!v8) | (!v1&!v2&!v3&!v5
    &v6&v7&!v8&v9) | (v2&v4&!v5&v6&!v7&v8&!v9));

hex[2] <= v0 ? ((!v1&v1&!v3&!v4&!v5&v6&v7&!v8&v9) | (!v1&v1&v3&v4&!v5&v6&!v7&!v8
    &!v9) | (v1&v1&!v3&!v4&!v5&!v6&!v7&!v8&v9) | (!v1&v1&!v3&v4&!v5&!v7
    &!v8&v9) | (v1&v1&!v3&!v4&v5&v6&v7&v8&v9) | (!v1&v1&!v3&v4&v5&!v6&!v7
    &v8&!v9) | (!v1&v1&!v3&v4&v5&!v6&v7&!v8&!v9) | (!v1&v1&!v3&v4&v5&v6
    &v7&!v8&v9) | (v1&!v1&!v3&v4&!v5&!v6&v7&v8&v9) | (v1&!v1&v3&v5&!v6&v7
    &!v8&!v9) | (v1&v1&!v4&!v5&v6&!v7&v8&!v9) | (v1&v3&v4&v5&v6&!v7&v8&!v9) | (
    !v1&v1&v3&v4&!v5&v7&v8&!v9) | (v1&!v3&!v4&!v5&v6&v7&v8&v9) | (v1&v1
    &v3&v4&v5&v6&!v8&!v9) | (!v1&v1&!v3&!v4&v5&!v6&!v7&!v8) | (v1&!v1&v3
    &v4&v6&!v7&v8&v9) | (v1&!v1&!v4&!v5&v6&!v7&!v8&v9) | (v1&v3&v4&!v5&v6
    &v7&v8&!v9) | (v1&!v1&!v3&v4&!v6&v7&v8&!v9) | (!v1&v1&!v3&v4&v6&v7&v8
    &!v9) | (!v1&!v3&v4&v5&v6&!v7&!v8&!v9) | (v1&v1&!v3&v4&v5&v6&!v7&v8) | (
    v1&!v1&!v3&v4&!v6&v7&!v8&v9) | (v1&!v1&!v3&v4&!v5&v6&!v7&v9) | (!v1
    &v1&v4&!v5&!v6&!v8&v9) | (v1&!v3&v4&!v5&v6&v7&!v8&v9) | (v1&v1&v3&!v4
    &v5&!v6&v7&!v8&v9) | (v1&!v1&v3&v4&v5&v6&v7&!v8&!v9) | (v1&!v1&!v3&!v4
    &!v5&!v6&!v7&v8&v9) | (v1&!v1&v3&!v4&!v6&v7&!v8&!v9) | (!v1&v1&v3&v5
    &!v6&!v7&v8&v9) | (v1&v3&!v4&!v5&v6&!v7&v8&v9) | (!v1&v1&!v3&!v4&!v5
    &!v6&v7&!v9) | (!v1&!v3&!v4&!v5&!v6&v7&v8&!v9) | (v1&!v1&!v3&!v4&v5
    &!v7&!v8&v9) | (v1&!v1&v3&v4&!v6&v7&v8&v9) | (v1&!v1&v3&v4&v5&v6&!v8
    &v9) | (!v1&v1&v3&v4&!v6&v7&!v8&v9) | (v1&v3&!v4&v5&v6&v7&!v8&!v9) | (
    !v1&!v1&!v3&v4&v6&!v7&!v8&!v9) | (!v1&!v1&!v4&v5&v6&v7&!v8&v9) | (v1
    &!v1&!v4&!v5&!v6&v7&v8&!v9) | (v1&v1&!v3&!v4&v5&v6&v7&!v9) | (v1&v1
    &!v3&v4&!v5&!v7&v8&!v9) | (v1&v1&!v4&v5&!v6&!v7&v8&v9) | (v1&v1&v3&v4
    &v5&v7&v8&v9) | (v1&!v1&v3&v4&!v5&v6&!v7&!v9) | (!v1&!v1&v3&!v5&v6&!v7
    &!v8&v9) | (v1&v3&v4&v5&!v6&!v7&!v8&!v9) | (v1&!v3&v4&v5&v6&v7&v8&v9) | (
    !v1&!v3&v4&v5&v6&!v7&!v8&!v9) | (!v1&v1&!v3&v4&!v5&v6&v7&!v9) | (!v1
    &v1&v3&!v4&v5&!v8&!v9) | (v1&!v1&!v3&v4&!v5&!v6&!v7&!v9) | (!v1&!v1
    &!v3&v4&v5&!v6&!v7&!v8) | (!v1&!v1&v3&v5&!v6&v8&!v9) | (v1&v3&!v4&v5
    &!v6&v8&v9) | (!v1&!v1&!v3&v4&!v5&v7&!v8&v9) | (v1&v1&!v3&v4&!v5&v6
    &!v8&!v9) | (!v1&!v4&v5&!v6&v7&!v8&!v9) | (!v1&!v1&v3&!v5&v6&v8&!v9) | (
    !v1&!v1&!v3&!v4&!v6&v8&v9) | (!v1&!v1&v3&!v5&v7&v8&v9) | (!v1&v3&!v4
    &!v5&!v6&!v7&v8) | (!v1&v1&!v3&!v4&v6&!v7&!v9) | (!v1&!v1&v3&v4&v5&v6
    &!v7) | (v1&!v3&!v4&v5&v6&!v8&!v9) | (v1&!v3&!v4&v6&v7&!v8&!v9) | (
    !v1&!v1&!v3&v5&v6&!v7&v8) | (!v1&!v1&!v3&!v4&!v5&!v6&!v8) | (!v1&!v1
    &!v3&v6&!v7&v8&v9) | (!v1&v1&v3&!v5&!v6&v7&!v8) | (!v1&v3&v4&!v5&!v6
    &v7&!v8) | (v1&v3&v4&!v5&!v6&!v7&v8) | (v1&!v1&!v3&v4&!v5&v8&!v9) | (
    !v1&!v1&!v3&!v6&!v7&!v8&v9) | (v1&v1&!v3&v5&!v6&v7&!v8) | (!v1&v1&!v3
    &v4&!v5&!v6&!v7) | (v1&v1&!v3&!v4&!v6&!v7&v8&!v9) | (v1&v1&v3&!v4&!v6
    &v8&v9) | (!v1&v3&v5&v6&v7&v8&!v9) | (!v1&!v1&v3&!v6&!v7&v8&!v9) | (
    !v1&!v1&v3&!v4&!v6&!v7&!v8) | (!v1&v1&!v3&!v4&!v5&v8&!v9) | (!v1&!v1
    &v3&!v4&!v5&!v7&!v8) | (v1&v1&v5&!v6&v7&v8&!v9) | (v1&!v3&!v4&!v5&!v6
    &v8&!v9) | (!v1&!v1&v4&v5&!v6&!v7&v9) | (v1&v1&!v3&v5&v7&!v8&!v9) | (
    !v1&v1&v4&!v5&!v6&v7&v9) | (v1&v1&v4&v5&!v6&!v7&!v8)) :
    ((v1&v2&!v3&!v5&v6&!v7&v8&v9) | (!v1&!v2&v3&v4&v6&v7&v8&!v9) | (v1
    &v2&!v3&!v4&v5&v6&!v7&v8&v9) | (v1&v2&v3&!v4&!v5&v6&!v7&!v8&!v9) | (
    v1&v2&!v3&!v4&!v5&!v6&v7&!v8&!v9) | (!v1&!v2&v3&!v4&!v5&!v6&v7&v8&!v9) | (
    !v1&v2&!v3&!v4&!v5&!v6&!v7&!v8&!v9) | (!v1&v2&v3&v4&v5&!v6&!v7&!v8&!v9) | (
    v1&!v2&v3&!v4&!v5&!v6&!v7&!v8&v9) | (!v1&!v2&v3&!v4&!v5&v6&v7&!v8&!v9) | (
    !v1&v2&v3&v4&!v5&!v6&!v7&v8&!v9) | (!v1&v2&!v3&!v4&!v5&!v6&!v7&v8&v9) | (
    !v1&v2&v3&!v4&!v5&!v6&!v7&!v8&!v9) | (v1&v2&v3&v4&v5&!v7&v8&!v9) | (
    v1&!v2&!v3&v4&!v5&v7&v8&!v9) | (v1&!v2&!v3&!v4&!v6&!v7&v8&!v9) | (!v1
    &!v2&!v3&v4&v6&!v7&v8&!v9) | (v1&!v2&v3&v4&v5&v6&!v7&v9) | (v1&!v2&!v3
    &!v4&!v6&v7&v8&v9) | (!v1&v2&!v3&!v4&v5&!v6&!v7&!v9) | (!v1&!v2&!v3
    &v4&!v5&!v7&!v8&!v9) | (!v1&v2&v3&!v4&v5&!v6&v8&!v9) | (!v1&v2&!v3&v4
    &v5&!v6&v7&!v9) | (!v1&v2&!v3&!v4&v5&v6&v7&v8) | (v1&!v2&!v4&!v5&v6
    &v7&!v8&v9) | (!v1&!v3&!v4&v5&v6&!v7&!v8&!v9) | (v1&v2&v3&!v5&!v6&v7
    &v8&v9) | (!v1&!v2&v3&!v4&!v5&!v6&v8&v9) | (!v1&v2&v3&v4&!v5&!v6&!v8
    &!v9) | (!v1&v2&v4&v5&v6&v7&!v8&v9) | (!v1&v2&v3&v4&v6&v7&!v8&!v9) | (
    !v1&v2&!v3&v4&v6&v7&!v8&v9) | (!v1&!v2&v3&v4&!v5&v6&!v8&v9) | (!v2&v3
    &!v4&v5&v6&v7&!v8&v9) | (!v1&!v2&v3&v5&v6&!v7&!v8&!v9) | (!v1&!v2&!v3
    &v5&!v6&v7&!v8&!v9) | (!v1&!v2&!v3&!v5&!v6&v7&!v8&v9) | (v1&v2&v3&!v4
    &v5&!v6&!v7&!v8&!v9) | (!v1&!v2&v3&v4&!v5&!v6&v7&!v8&!v9) | (v1&v2&!v4
    &!v5&v6&v7&v8&!v9) | (v1&!v2&!v3&v4&!v5&v6&v7&!v9) | (v1&!v2&!v3&v4
    &v5&!v6&v8&v9) | (v1&!v2&!v4&v5&v6&v7&v8&v9) | (v1&!v2&!v3&v4&!v5&!v6
    &!v7&v9) | (v1&!v2&v3&v4&!v5&!v7&!v8&!v9) | (v2&v3&v4&v5&v6&v7&v8&!v9) | (
    v1&!v2&!v3&v5&!v6&v7&v8&!v9) | (!v1&!v2&!v3&!v4&v6&v7&v8&!v9) | (!v1
    &v2&v3&v4&!v6&!v7&v8&v9) | (!v2&!v3&!v4&!v5&v6&!v7&!v8&!v9) | (!v1&!v2
    &v3&v4&v5&!v6&v7&v8) | (!v1&!v3&v4&v5&v6&!v7&!v8&v9) | (v1&v2&!v4&!v5
    &v6&!v7&v8&v9) | (!v1&v3&!v4&!v5&v6&!v7&!v8&v9) | (v1&v2&!v3&!v4&!v6
    &v7&v8&!v9) | (v1&!v2&v3&!v4&v5&v6&!v7&!v9) | (v1&v2&!v3&!v4&v5&v6&v7
    &!v9) | (v1&v2&!v3&v4&!v5&!v6&!v8&!v9) | (!v1&v2&!v3&v4&v5&!v6&!v7&v8) | (
    v1&!v2&v3&v5&!v6&!v7&v8&v9) | (!v1&!v2&!v3&!v4&!v5&v6&!v7&v9) | (!v1
    &!v2&!v3&v5&v6&v7&v8&!v9) | (!v1&!v2&!v3&v4&v5&!v6&!v7&!v8) | (!v1&v2
    &v3&v4&!v6&!v7&!v8&v9) | (v1&v2&!v3&!v4&!v5&!v7&v9) | (v1&v3&!v4&!v5
    &!v6&v8&!v9) | (!v2&!v3&!v4&!v5&!v7&v8&v9) | (v1&!v2&!v3&v4&!v7&!v8
    &v9) | (!v1&v3&!v4&v5&!v7&v8&v9) | (!v1&v2&!v3&v4&!v6&v8&v9) | (v1&!v2
    &v3&v4&!v6&!v8&!v9) | (v1&v2&!v4&v5&!v6&!v8&v9) | (!v1&v2&v3&!v4&v6
    &!v7&v8) | (v1&v2&v3&!v4&!v6&v7&v9) | (!v1&v3&v4&v5&v6&v7&v8) | (!v2
    &!v3&!v4&v5&!v6&v7&v9) | (!v2&!v3&v4&v5&v6&v7&!v8) | (v2&!v3&v5&v6&!v7
    &!v8&!v9) | (v1&!v2&v3&v5&v7&!v8&!v9) | (v1&v2&!v3&v5&v7&!v8&v9) | (
    v1&!v2&!v3&v5&!v6&!v7&!v8) | (!v1&v2&v3&!v5&v6&!v7&v9) | (v2&v3&!v4
    &v5&!v6&v7&!v8) | (v2&v3&!v5&!v6&!v7&!v8&v9) | (v1&!v3&v4&!v5&v6&v7
    &v8&!v9) | (!v1&!v2&v4&v5&v6&!v7&!v8&v9) | (v2&!v3&!v4&v5&v6&v7&!v8
    &v9) | (v1&v3&v4&v5&v6&!v7&v8) | (!v1&v3&v4&!v5&!v6&!v7&v9) | (v2&v3
    &!v4&v5&v7&!v8&!v9) | (v1&v2&v3&!v4&v5&v8&v9) | (!v1&v2&!v3&!v4&!v5
    &v7&!v9) | (v1&v2&!v4&v5&v7&!v8&v9) | (v1&!v2&!v3&!v6&!v7&!v8&v9));

hex[1] <= v0 ? ((!v1&v1&v3&v4&v5&v6&!v7&!v8&v9) | (v1&v1&!v3&!v4&v5&v6&v7&v8&v9) | (
    !v1&v1&!v3&v4&v5&!v6&!v7&v8&!v9) | (!v1&v1&!v3&v4&v5&!v6&v7&!v8&!v9) | (
    !v1&v3&!v4&v5&!v6&!v7&!v8&!v9) | (v1&v1&!v3&v4&v5&!v6&v7&!v8&v9) | (
    v1&!v1&v3&!v4&!v5&v6&!v7&!v9) | (!v1&v1&!v3&!v4&v5&!v6&v7&v8) | (!v1
    &!v3&!v4&v5&v6&v7&!v8&v9) | (v1&v1&!v3&!v4&v5&!v7&!v8&!v9) | (!v1&v3
    &v4&!v5&!v6&v7&v8&v9) | (v1&!v1&!v3&v4&v5&!v7&v8&!v9) | (!v1&v1&!v3
    &v4&v5&v7&v8&v9) | (!v1&v1&v4&!v5&v6&v7&v8&!v9) | (v1&v1&!v3&!v4&v6
    &!v7&!v8&v9) | (!v1&!v1&!v3&!v5&!v6&!v7&v8&v9) | (!v1&v3&v4&!v5&v6&v7
    &!v8&v9) | (v1&v1&v4&!v5&v6&v7&v8&v9) | (v1&!v3&v4&!v5&v6&v7&!v8&!v9) | (
    v1&v1&!v3&v4&!v6&!v7&!v8&!v9) | (v1&v1&v3&!v4&v5&!v6&v7&!v8&v9) | (
    v1&!v1&v3&v4&v5&v6&v7&!v8&!v9) | (v1&!v1&!v3&!v4&!v5&!v6&!v7&v8&v9) | (
    v1&!v1&v3&!v4&!v6&v7&!v8&!v9) | (!v1&v1&v3&v5&!v6&!v7&v8&v9) | (v1&v3
    &!v4&!v5&v6&!v7&v8&v9) | (!v1&v1&!v3&!v4&!v5&!v6&v7&!v9) | (!v1&!v3
    &!v4&!v5&!v6&v7&v8&!v9) | (v1&!v1&!v3&!v4&v5&!v7&!v8&v9) | (v1&!v1&v3
    &v4&!v6&v7&v8&v9) | (v1&!v1&v3&!v4&v6&v7&v8&!v9) | (v1&!v1&v3&v4&v5
    &v6&!v8&v9) | (!v1&v1&v3&v4&!v6&v7&!v8&v9) | (!v1&!v1&v3&v5&v6&!v7&!v8
    &!v9) | (v1&!v1&!v4&v5&v6&v7&!v8&v9) | (v1&!v1&v3&v5&v6&!v7&v8&v9) | (
    !v1&!v1&!v3&v4&v6&!v7&!v8&!v9) | (v1&v1&!v3&v4&!v5&!v7&v8&!v9) | (!v1
    &!v1&!v3&v4&v5&v6&v8&!v9) | (v1&v3&v4&v5&!v6&!v7&!v8&v9) | (v1&v1&!v3
    &!v4&!v5&!v7&v8&v9) | (!v1&v1&v3&v4&!v5&!v6&!v8&!v9) | (v1&!v3&!v4&!v5
    &!v6&v7&!v8&v9) | (v1&!v3&v4&v5&v6&!v7&v8&v9) | (v1&!v1&v3&v4&!v5&v6
    &v7&!v8) | (v1&!v3&v4&v5&v6&v7&!v8&!v9) | (!v1&!v3&v4&!v5&v6&v7&!v8
    &!v9) | (v1&v1&v3&v5&!v6&v8&!v9) | (v1&v1&v3&!v4&!v6&v7&v8) | (v1&v3
    &v5&!v6&v7&v8&!v9) | (v1&!v1&!v3&!v4&!v6&v8&!v9) | (!v1&!v1&v3&!v4&!v5
    &!v6&!v8) | (!v1&!v1&!v4&v5&v6&!v7&!v8) | (!v1&!v1&v3&v4&!v5&v8&!v9) | (
    !v1&v3&v4&v5&!v6&v7&v9) | (v1&!v3&v4&!v5&v6&!v7&!v8&v9) | (!v1&!v1&!v3
    &v4&v5&v7&!v9) | (v1&v3&!v4&!v5&v7&!v8&v9) | (!v1&!v3&!v4&!v5&!v7&v8
    &v9) | (v1&v3&!v4&!v5&!v6&!v7&!v8) | (!v1&!v3&v5&v6&!v7&v8&v9) | (v1
    &!v1&v4&v5&!v6&v7&v9) | (v1&v1&v3&v4&v5&v6&v7) | (!v1&!v1&!v5&v6&v7
    &v8&v9) | (v1&v3&!v5&v6&!v7&v8&!v9) | (v1&!v1&v4&v6&v7&v8&!v9) | (v1
    &!v1&v4&v5&v6&!v7&v9) | (v1&v3&v4&!v5&!v6&!v8&!v9) | (v1&!v1&!v3&!v6
    &v7&!v8&!v9) | (!v1&!v1&!v3&!v5&v7&!v8&v9) | (!v1&!v3&v4&v5&!v6&!v7
    &!v8) | (!v1&v4&!v5&!v6&!v7&!v8&v9) | (v1&v1&!v3&v4&!v5&!v6&v8) | (
    v1&v1&!v3&!v4&!v6&!v7&v8&!v9) | (v1&v1&v3&!v4&!v6&v8&v9) | (!v1&v3&v5
    &v6&v7&v8&!v9) | (!v1&!v1&v3&!v6&!v7&v8&!v9) | (!v1&!v1&v3&!v4&!v6&!v7
    &!v8) | (!v1&v1&!v3&!v4&!v5&v8&!v9) | (!v1&!v1&v3&!v4&!v5&!v7&!v8) | (
    v1&v1&v5&!v6&v7&v8&!v9) | (!v1&!v1&v3&v4&v5&!v7&v8) | (!v1&!v3&!v4&v5
    &v7&!v8) | (v3&v4&!v5&!v7&v8&!v9) | (!v1&!v5&v6&!v7&!v8&!v9)) :
    ((v1&!v2&v3&!v4&v5&!v7&!v8&!v9) | (!v1&v2&!v3&!v4&!v5&v6&v7&v9) | (
    v1&v2&!v3&!v4&v5&v6&!v7&v8&v9) | (v1&v2&v3&!v4&!v5&v6&!v7&!v8&!v9) | (
    v1&v2&!v3&!v4&!v5&!v6&v7&!v8&!v9) | (!v1&!v2&v3&!v4&!v5&!v6&v7&v8&!v9) | (
    !v1&v2&!v3&!v4&!v5&!v6&!v7&!v8&!v9) | (!v1&v2&v3&v4&v5&!v6&!v7&!v8&!v9) | (
    v1&!v2&v3&!v4&!v5&!v6&!v7&!v8&v9) | (!v1&!v2&v3&!v4&!v5&v6&v7&!v8&!v9) | (
    v1&v2&!v4&v5&!v6&v7&v8&!v9) | (!v1&!v2&!v3&v4&!v5&!v7&v8&!v9) | (v1
    &v2&!v3&v4&v6&!v7&!v8&!v9) | (v1&!v2&!v3&!v4&!v6&v7&v8&!v9) | (!v1&v2
    &v4&!v5&v6&!v7&v8&v9) | (v1&!v2&v3&v4&v5&v7&v8&v9) | (v1&!v2&v3&!v4
    &v5&!v6&!v7&!v9) | (!v1&v2&!v3&v4&v5&v6&!v7&v8) | (v1&v3&v4&!v5&!v6
    &!v7&!v8&!v9) | (!v2&!v3&v4&!v5&v6&v7&v8&v9) | (!v1&!v2&!v3&!v4&v5&!v6
    &!v7&!v9) | (v1&!v2&v3&!v5&v6&v7&v8&!v9) | (v1&v2&!v3&v4&v5&!v6&v7&!v8) | (
    !v1&v2&v4&!v5&!v6&!v7&!v8&v9) | (!v1&v2&!v4&!v5&v6&v7&!v8&!v9) | (!v1
    &v2&v3&v5&!v6&!v7&v8&!v9) | (!v1&!v2&!v3&!v4&!v6&v7&v8&v9) | (v1&!v2
    &!v3&!v4&v5&!v6&v7&!v8) | (!v2&v3&v4&v5&!v6&!v7&!v8&v9) | (v1&!v2&v3
    &!v5&!v6&v7&v8&v9) | (v1&v2&v3&!v4&v5&!v6&!v7&!v8&!v9) | (!v1&!v2&v3
    &v4&!v5&!v6&v7&!v8&!v9) | (v1&v2&!v4&!v5&v6&v7&v8&!v9) | (v1&!v2&!v3
    &v4&!v5&v6&v7&!v9) | (v1&!v2&!v3&v4&v5&!v6&v8&v9) | (v1&!v2&!v4&v5&v6
    &v7&v8&v9) | (v1&!v2&!v3&v4&!v5&!v6&!v7&v9) | (v1&!v2&v3&v4&!v5&!v7
    &!v8&!v9) | (v2&v3&v4&v5&v6&v7&v8&!v9) | (v1&!v2&!v3&v5&!v6&v7&v8&!v9) | (
    !v1&!v2&!v3&!v4&v6&v7&v8&!v9) | (!v1&v2&v3&v4&!v6&!v7&v8&v9) | (!v2
    &!v3&!v4&!v5&v6&!v7&!v8&!v9) | (!v1&!v2&v3&v4&v5&!v6&v7&v8) | (!v1&!v3
    &v4&v5&v6&!v7&!v8&v9) | (v1&!v2&!v4&v5&v6&!v7&v8&v9) | (v1&v2&v3&!v4
    &!v5&v6&!v7&v8) | (!v1&v3&!v4&!v5&v6&!v7&!v8&v9) | (!v1&v2&v4&!v5&!v6
    &v7&v8&v9) | (!v1&!v2&v4&v5&!v6&!v7&!v8&!v9) | (!v1&v3&!v4&!v5&!v6&!v7
    &v8&v9) | (!v1&!v2&!v3&v4&!v5&v6&!v8&!v9) | (!v1&v2&v3&v4&!v5&v6&!v8
    &!v9) | (!v1&v2&v3&!v4&v5&v6&!v7&!v8) | (v2&v3&!v4&!v5&!v6&v7&!v8&v9) | (
    v1&v4&v5&v6&!v7&v8&!v9) | (!v2&!v4&!v5&v6&!v7&v8&!v9) | (v1&!v3&v4&!v5
    &v6&v8&v9) | (!v1&v2&v4&!v5&v7&v8&!v9) | (v1&v2&!v3&!v4&v5&!v6&v8) | (
    !v1&!v2&!v4&v6&!v7&v8&!v9) | (v1&v2&v3&!v4&v6&v7&v8) | (!v1&!v3&!v4
    &!v5&v6&!v7&!v9) | (!v2&v3&v4&!v5&!v6&v8&v9) | (v1&!v2&!v3&!v5&!v6&!v7
    &v8) | (v2&v3&v4&!v5&!v6&v7&v8) | (v1&v2&v4&!v6&v7&!v8&v9) | (v1&v3
    &v4&v6&v7&!v8&v9) | (!v1&!v3&v5&!v6&v7&v8&!v9) | (!v1&!v2&!v4&!v5&!v6
    &!v7&!v8) | (!v1&!v2&!v3&!v4&v5&!v8&v9) | (!v1&v2&!v3&!v4&!v5&v6&!v8) | (
    v1&!v2&!v3&!v5&v7&!v8&v9) | (!v2&!v3&v5&v6&!v7&!v8&v9) | (!v1&!v2&v3
    &v5&!v6&v8&v9) | (v2&v3&!v5&v6&!v7&!v8&v9) | (!v1&!v2&v3&v5&v7&!v8&!v9) | (
    v2&v3&v5&!v6&v7&!v8&v9) | (!v2&v3&!v5&v6&v7&!v8&v9) | (v1&!v3&v4&!v5
    &v6&v7&v8&!v9) | (!v1&!v2&v4&v5&v6&!v7&!v8&v9) | (v2&!v3&!v4&v5&v6&v7
    &!v8&v9) | (v1&v3&v4&v5&v6&!v7&v8) | (!v1&v3&v4&!v5&!v6&!v7&v9) | (
    v2&v3&!v4&v5&v7&!v8&!v9) | (v1&v2&!v3&v5&v6&!v7&!v9) | (!v2&!v3&!v4
    &v5&v6&v7&!v9) | (v1&!v3&v5&!v6&!v7&v8&v9) | (v1&v2&v3&v4&v5&v6) | (
    v3&!v4&v5&v6&v7&!v9));

hex[0] <= v0 ? ((!v1&!v1&!v3&!v5&!v6&v7&!v8&!v9) | (v1&!v1&v3&v4&v5&v6&v7&v8&v9) | (
    !v1&v1&!v3&!v4&!v5&!v6&!v7&!v8&!v9) | (v1&!v1&!v3&!v4&!v5&!v6&v7&!v8
    &v9) | (v1&v1&v3&v4&!v5&!v6&v7&v8&v9) | (!v1&!v1&!v3&v4&!v5&v6&!v7&v8
    &!v9) | (v1&!v1&!v3&v4&!v5&v6&v7&v8&v9) | (!v1&v1&!v3&v4&!v5&v6&v7&v8
    &v9) | (v1&!v1&!v3&v4&!v5&v6&!v7&!v8&!v9) | (v1&v1&!v3&v4&v5&!v6&v7
    &!v8&v9) | (!v1&v1&!v3&v4&v5&v6&v7&!v8&v9) | (v1&!v1&!v3&v4&!v5&!v6
    &v7&v8&v9) | (!v1&v3&!v4&v5&!v6&v7&v8&!v9) | (v1&!v1&!v4&v5&v6&v7&v8
    &!v9) | (!v1&v3&!v4&!v5&v6&v7&!v8&!v9) | (v1&v3&!v4&!v5&!v6&v7&!v8&!v9) | (
    !v1&!v1&!v3&!v4&v5&v6&v7) | (!v1&!v1&v3&!v5&!v6&v7&!v8&v9) | (!v1&!v3
    &!v4&!v5&v6&!v7&!v8&!v9) | (v1&v1&v3&v4&!v5&v7&v8&!v9) | (!v1&!v1&v3
    &v4&!v5&v6&v7&v8) | (!v1&!v1&!v3&v4&!v5&!v6&v7&!v9) | (v1&v1&v3&!v4
    &v5&!v6&v7&!v8&v9) | (v1&v1&v3&v4&!v5&!v7&!v8&v9) | (v1&!v1&v3&v4&v5
    &v6&v7&!v8&!v9) | (v1&!v1&!v3&!v4&!v5&!v6&!v7&v8&v9) | (!v1&!v3&v4&!v5
    &!v6&!v7&!v8&v9) | (!v1&!v1&!v3&!v4&v5&!v6&v8&!v9) | (!v1&!v3&!v4&v5
    &!v6&!v7&!v8&!v9) | (v1&!v1&!v3&!v4&v6&!v7&v8&v9) | (!v1&v1&v3&!v5&!v6
    &!v7&v8&v9) | (!v1&v1&!v3&v5&!v6&!v7&v8&v9) | (v1&v1&!v3&!v4&v6&v7&!v8
    &v9) | (v1&!v1&v3&!v4&v6&v7&v8&!v9) | (v1&v3&v4&!v5&v6&v7&!v8&v9) | (
    !v1&!v1&v3&v5&v6&!v7&!v8&!v9) | (v1&!v1&!v4&v5&v6&v7&!v8&v9) | (v1&!v1
    &v3&v5&v6&!v7&v8&v9) | (v1&v3&!v4&v5&v6&v7&!v8&!v9) | (!v1&!v1&!v4&v5
    &v6&v7&!v8&v9) | (v1&!v1&!v4&!v5&!v6&v7&v8&!v9) | (v1&v1&!v3&!v4&v5
    &v6&v7&!v9) | (v1&v1&!v4&v5&!v6&!v7&v8&v9) | (!v1&!v1&!v3&v4&v5&v6&v8
    &!v9) | (v1&v1&v3&v4&v5&v7&v8&v9) | (v1&v3&v4&v5&!v6&!v7&!v8&v9) | (
    v1&v1&!v3&!v4&!v5&!v7&v8&v9) | (!v1&v1&v3&v4&!v5&!v6&!v8&!v9) | (v1
    &!v1&v3&v4&!v5&v6&!v7&!v9) | (!v1&!v1&v3&!v5&v6&!v7&!v8&v9) | (v1&!v3
    &!v4&!v5&!v6&v7&!v8&v9) | (v1&!v3&v4&v5&v6&!v7&v8&v9) | (v1&v3&v4&v5
    &!v6&!v7&!v8&!v9) | (v1&!v1&v3&v4&!v5&v6&v7&!v8) | (v1&!v3&v4&v5&v6
    &v7&v8&v9) | (v1&!v3&v4&v5&v6&v7&!v8&!v9) | (!v1&!v3&v4&v5&v6&!v7&!v8
    &!v9) | (!v1&v1&!v3&v4&!v5&v6&v7&!v9) | (v1&!v1&!v3&v4&!v5&!v6&!v7&!v9) | (
    !v1&!v1&!v3&v4&v5&!v6&!v7&!v8) | (!v1&!v3&v4&!v5&v6&v7&!v8&!v9) | (
    !v1&!v1&!v3&v4&!v5&v7&!v8&v9) | (v1&v1&!v3&v4&!v5&v6&!v8&!v9) | (v1
    &!v3&v4&!v5&v6&!v7&!v8&v9) | (!v1&v3&!v4&v5&!v6&v8&v9) | (!v1&!v3&!v4
    &v5&v6&v8&v9) | (!v1&v1&v3&!v4&!v5&!v7&v9) | (!v1&v1&v3&!v4&!v5&v7&v8) | (
    !v1&v3&!v4&!v6&!v7&!v8&!v9) | (!v1&!v3&!v4&v5&v7&!v8&v9) | (v1&v1&v3
    &!v4&v5&!v7&!v8) | (v1&!v1&!v4&v5&!v6&v7&!v8) | (v1&!v1&!v4&!v5&v6&v7
    &v9) | (!v1&!v1&!v3&!v4&v6&v7&v8) | (v1&!v1&!v3&!v4&v5&!v6&!v7) | (
    !v1&v1&!v4&!v5&!v6&!v7&v9) | (v1&!v1&v3&!v4&!v5&!v7&!v8) | (v1&v1&v5
    &v6&!v7&v8&!v9) | (!v1&!v1&v3&!v5&!v6&!v7&v8) | (v1&!v4&!v5&!v6&!v7
    &!v8&!v9) | (v1&!v1&v3&v4&!v7&v8&v9) | (!v1&v3&v4&!v5&!v6&!v7&!v9) | (
    v1&!v1&!v4&!v5&v6&v7&!v8) | (v1&!v1&!v3&!v6&!v7&v8&!v9) | (!v1&!v1&v4
    &v5&!v6&v7&!v8) | (v1&!v3&v5&v6&!v7&!v8&!v9) | (v1&v1&v4&v5&!v6&!v8
    &!v9) | (v1&!v3&v4&v5&!v6&v8&!v9) | (!v1&v1&!v3&!v5&!v7&v8&!v9) | (
    v1&v1&!v3&!v6&!v7&v8&v9) | (!v1&v1&v4&!v5&v7&!v8&!v9) | (!v1&v1&!v3
    &!v5&v6&!v8&!v9) | (v1&!v3&!v5&!v6&v7&v8&v9) | (v1&v4&!v5&v6&!v7&v8
    &!v9) | (v1&!v1&!v3&!v5&v6&!v7&v8) | (v1&v1&!v3&!v4&!v6&!v7&v8&!v9) | (
    v1&v1&!v3&v4&!v5&v6&v7) | (!v1&v1&v3&v4&v5&v6&v7) | (!v1&!v1&v3&v4&v5
    &!v7&v8) | (v1&!v3&!v4&!v5&!v6&v8&!v9) | (!v1&!v1&v4&v5&!v6&!v7&v9) | (
    v1&v1&!v3&v5&v7&!v8&!v9) | (!v1&v1&v4&!v5&!v6&v7&v9) | (v1&v1&v4&v5
    &!v6&!v7&!v8) | (v1&!v4&v5&v6&!v7&v9) | (!v1&v1&v3&v4&v5&v9) | (v1&v3
    &!v4&v6&v7&!v8) | (v1&v3&v5&v6&v7&v9) | (!v1&!v1&!v3&v5&v7&v9) | (!v1
    &v3&v4&v5&v6&!v7) | (!v1&!v1&v4&v5&!v8&v9) | (v1&!v4&!v5&!v6&!v7&v8) | (
    !v1&v3&v4&v6&!v7&!v8) | (v1&!v3&v6&!v7&v8&!v9)):
    ((v1&!v2&v3&v4&!v5&!v6&!v7&v8&!v9) | (v1&v2&!v3&!v4&v5&v6&v7&v8&v9) | (
    v1&v2&!v3&!v4&!v5&v6&!v7&!v8&!v9) | (!v1&!v2&!v3&v4&v5&v6&!v7&!v8&!v9) | (
    v1&!v2&v3&!v4&!v5&v6&!v7&!v8&v9) | (!v1&v2&v3&!v4&!v5&v6&!v7&!v8&!v9) | (
    !v1&v2&v3&v4&!v5&!v6&!v7&v8&!v9) | (!v1&v2&!v3&!v4&!v5&!v6&!v7&v8&v9) | (
    !v1&v2&v3&!v4&!v5&!v6&!v7&!v8&!v9) | (v1&v3&v4&!v5&v6&!v7&v8&v9) | (
    v1&v2&v3&v4&v5&!v6&v7&!v9) | (v1&!v2&v3&v4&v5&v6&v7&v8) | (v1&!v2&v3
    &!v4&!v6&v7&v8&!v9) | (v1&!v2&v3&v4&!v5&!v6&v7&v9) | (v2&!v3&!v4&v5
    &!v6&!v7&!v8&!v9) | (v1&v3&v4&!v5&!v6&v7&!v8&!v9) | (v1&!v2&v3&v5&v6
    &v7&v8&!v9) | (!v1&!v2&v3&!v4&v5&v6&v8&v9) | (!v1&v2&!v3&v4&!v6&v7&!v8
    &!v9) | (v1&!v2&v3&!v5&!v6&!v7&!v8&!v9) | (!v1&!v2&!v4&!v5&!v6&v7&!v8
    &v9) | (!v1&v2&!v3&v5&v6&v7&!v8&!v9) | (!v1&!v2&v3&v5&v6&v7&!v8&!v9) | (
    !v1&v2&!v3&v5&!v6&v7&!v8&v9) | (v1&v2&v3&!v4&v5&!v6&!v7&!v8&!v9) | (
    !v1&!v2&v3&v4&!v5&!v6&v7&!v8&!v9) | (v1&v2&!v3&v4&!v5&!v6&!v7&v9) | (
    !v1&v2&!v4&!v5&!v6&!v7&v8&!v9) | (v1&!v3&v4&!v5&!v6&v7&v8&v9) | (!v1
    &!v2&v4&v5&v6&!v7&v8&v9) | (!v1&v2&v3&v4&v5&v6&!v7&!v9) | (!v1&!v2&!v3
    &v4&v6&!v7&v8&v9) | (!v1&!v3&v4&v5&v6&v7&v8&v9) | (v1&v3&!v4&!v5&v6
    &v7&!v8&!v9) | (!v1&!v2&!v3&!v4&v6&v7&v8&v9) | (v1&v2&v3&!v4&!v5&v6
    &v7&!v8) | (!v1&v2&!v4&v5&!v6&!v7&!v8&v9) | (!v1&!v2&v3&!v4&v5&!v6&!v7
    &!v8) | (v1&!v2&!v4&v5&v6&!v7&v8&v9) | (!v1&!v2&!v3&!v5&v6&v7&!v8&v9) | (
    v1&v2&v3&!v4&!v5&v6&!v7&v8) | (v1&v2&!v4&!v5&v6&!v7&v8&v9) | (v1&v2
    &!v3&!v4&!v6&v7&v8&!v9) | (v1&!v2&v3&!v4&v5&v6&!v7&!v9) | (v1&v2&!v3
    &!v4&v5&v6&v7&!v9) | (!v1&v2&v4&!v5&!v6&v7&v8&v9) | (v1&v2&!v3&v4&!v5
    &!v6&!v8&!v9) | (!v1&v2&!v3&v4&v5&!v6&!v7&v8) | (!v1&!v2&v4&v5&!v6&!v7
    &!v8&!v9) | (!v1&v3&!v4&!v5&!v6&!v7&v8&v9) | (!v1&!v2&!v3&v4&!v5&v6
    &!v8&!v9) | (!v1&v2&v3&v4&!v5&v6&!v8&!v9) | (v1&!v2&v3&v5&!v6&!v7&v8
    &v9) | (!v1&!v2&!v3&!v4&!v5&v6&!v7&v9) | (!v1&v2&v3&!v4&v5&v6&!v7&!v8) | (
    !v1&!v2&!v3&v5&v6&v7&v8&!v9) | (!v1&!v2&!v3&v4&v5&!v6&!v7&!v8) | (v2
    &v3&!v4&!v5&!v6&v7&!v8&v9) | (!v1&v2&v3&v4&!v6&!v7&!v8&v9) | (v1&!v3
    &v4&v5&v6&!v7&v8) | (v1&!v2&!v3&v4&!v5&v6&!v9) | (v1&v2&v3&v4&!v5&v8
    &v9) | (v2&v3&v4&v5&!v7&v8&v9) | (v1&v2&!v3&!v6&!v7&v8&!v9) | (v1&!v2
    &v3&v4&v6&v7&!v9) | (v1&!v2&v3&!v4&v5&!v7&v9) | (v1&v2&!v3&v4&v6&v7
    &v9) | (!v1&!v3&v4&v5&!v6&!v7&!v9) | (!v1&!v2&v4&!v5&!v7&!v8&!v9) | (
    !v1&!v2&!v3&v4&!v5&v7&v8) | (v1&v4&!v5&v6&v7&!v8&v9) | (!v1&!v2&!v3
    &!v4&!v6&!v7&!v9) | (!v2&!v3&!v4&!v5&!v6&v7&!v9) | (!v1&v2&!v3&!v4&v6
    &v8&v9) | (v1&v3&v4&v5&!v6&!v7&!v8) | (!v1&v3&v4&!v5&v6&v7&v8) | (v2
    &!v3&v4&!v5&v6&!v8&v9) | (v3&!v4&v5&!v6&v7&v8&v9) | (v2&v3&v4&!v5&v6
    &!v7&!v8) | (!v1&v4&v5&!v6&v7&!v8&!v9) | (!v1&v2&!v3&!v5&v6&!v7&v8) | (
    v1&v3&!v4&!v5&!v6&!v8&v9) | (v1&v2&!v3&!v5&!v6&v7&v9) | (v1&v2&v3&v5
    &v6&!v8&!v9) | (!v1&v2&!v5&v6&v7&v8&v9) | (v1&v2&!v3&!v5&v6&v7&!v8) | (
    v1&!v2&!v3&v5&v6&v7&!v8) | (!v1&v2&v3&!v6&v7&v8&v9) | (!v1&!v2&!v3&v6
    &!v7&!v8&v9) | (v2&v3&v5&v6&v7&!v8&v9) | (!v1&!v2&v3&!v5&!v6&!v8&v9) | (
    v1&!v3&v4&!v5&v6&v7&v8&!v9) | (!v1&!v2&v4&v5&v6&!v7&!v8&v9) | (v2&!v3
    &!v4&v5&v6&v7&!v8&v9) | (v1&v2&!v3&v5&v6&!v7&!v9) | (v1&v2&v3&!v4&v5
    &v8&v9) | (!v2&!v3&!v4&v5&v6&v7&!v9) | (v1&!v3&v5&!v6&!v7&v8&v9) | (
    !v1&v2&!v3&!v4&!v5&v7&!v9) | (v1&v2&!v4&v5&v7&!v8&v9) | (v1&!v2&!v3
    &!v6&!v7&!v8&v9) | (v1&v2&v4&v5&!v7&v9) | (v1&v2&!v3&v4&v5&v8) | (!v3
    &!v4&v6&!v7&v8&!v9) | (!v2&!v3&!v4&v6&v8&!v9) | (v2&v3&!v4&v5&!v6&v8));

	end

	decoder decoder(.hex(hex), .segments(io_out));

endmodule

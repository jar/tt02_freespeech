module jar_pi
(
	input  [7:0] io_in,
	output [7:0] io_out
);
	wire       clk      = io_in[0];
	wire       reset    = io_in[1];
	wire       stream   = io_in[2];
	wire [4:0] io_index = io_in[7:3];

	reg [9:0] index;
	reg [7:0] led_out;
	reg [3:0] code;
	assign io_out[7:0] = led_out;

	always @(posedge clk) begin
		if (reset) begin
			index <= {io_index, index[9:5]};
		end
		else if (stream) begin
			index <= index + 1;

			case(index)
				   0: code <= 3;
				   1: code <= 10;
				   2: code <= 1;
				   3: code <= 4;
				   4: code <= 1;
				   5: code <= 5;
				   6: code <= 9;
				   7: code <= 2;
				   8: code <= 6;
				   9: code <= 5;
				  10: code <= 3;
				  11: code <= 5;
				  12: code <= 8;
				  13: code <= 9;
				  14: code <= 7;
				  15: code <= 9;
				  16: code <= 3;
				  17: code <= 2;
				  18: code <= 3;
				  19: code <= 8;
				  20: code <= 4;
				  21: code <= 6;
				  22: code <= 2;
				  23: code <= 6;
				  24: code <= 4;
				  25: code <= 3;
				  26: code <= 3;
				  27: code <= 8;
				  28: code <= 3;
				  29: code <= 2;
				  30: code <= 7;
				  31: code <= 9;
				  32: code <= 5;
				  33: code <= 0;
				  34: code <= 2;
				  35: code <= 8;
				  36: code <= 8;
				  37: code <= 4;
				  38: code <= 1;
				  39: code <= 9;
				  40: code <= 7;
				  41: code <= 1;
				  42: code <= 6;
				  43: code <= 9;
				  44: code <= 3;
				  45: code <= 9;
				  46: code <= 9;
				  47: code <= 3;
				  48: code <= 7;
				  49: code <= 5;
				  50: code <= 1;
				  51: code <= 0;
				  52: code <= 5;
				  53: code <= 8;
				  54: code <= 2;
				  55: code <= 0;
				  56: code <= 9;
				  57: code <= 7;
				  58: code <= 4;
				  59: code <= 9;
				  60: code <= 4;
				  61: code <= 4;
				  62: code <= 5;
				  63: code <= 9;
				  64: code <= 2;
				  65: code <= 3;
				  66: code <= 0;
				  67: code <= 7;
				  68: code <= 8;
				  69: code <= 1;
				  70: code <= 6;
				  71: code <= 4;
				  72: code <= 0;
				  73: code <= 6;
				  74: code <= 2;
				  75: code <= 8;
				  76: code <= 6;
				  77: code <= 2;
				  78: code <= 0;
				  79: code <= 8;
				  80: code <= 9;
				  81: code <= 9;
				  82: code <= 8;
				  83: code <= 6;
				  84: code <= 2;
				  85: code <= 8;
				  86: code <= 0;
				  87: code <= 3;
				  88: code <= 4;
				  89: code <= 8;
				  90: code <= 2;
				  91: code <= 5;
				  92: code <= 3;
				  93: code <= 4;
				  94: code <= 2;
				  95: code <= 1;
				  96: code <= 1;
				  97: code <= 7;
				  98: code <= 0;
				  99: code <= 6;
				 100: code <= 7;
				 101: code <= 9;
				 102: code <= 8;
				 103: code <= 2;
				 104: code <= 1;
				 105: code <= 4;
				 106: code <= 8;
				 107: code <= 0;
				 108: code <= 8;
				 109: code <= 6;
				 110: code <= 5;
				 111: code <= 1;
				 112: code <= 3;
				 113: code <= 2;
				 114: code <= 8;
				 115: code <= 2;
				 116: code <= 3;
				 117: code <= 0;
				 118: code <= 6;
				 119: code <= 6;
				 120: code <= 4;
				 121: code <= 7;
				 122: code <= 0;
				 123: code <= 9;
				 124: code <= 3;
				 125: code <= 8;
				 126: code <= 4;
				 127: code <= 4;
				 128: code <= 6;
				 129: code <= 0;
				 130: code <= 9;
				 131: code <= 5;
				 132: code <= 5;
				 133: code <= 0;
				 134: code <= 5;
				 135: code <= 8;
				 136: code <= 2;
				 137: code <= 2;
				 138: code <= 3;
				 139: code <= 1;
				 140: code <= 7;
				 141: code <= 2;
				 142: code <= 5;
				 143: code <= 3;
				 144: code <= 5;
				 145: code <= 9;
				 146: code <= 4;
				 147: code <= 0;
				 148: code <= 8;
				 149: code <= 1;
				 150: code <= 2;
				 151: code <= 8;
				 152: code <= 4;
				 153: code <= 8;
				 154: code <= 1;
				 155: code <= 1;
				 156: code <= 1;
				 157: code <= 7;
				 158: code <= 4;
				 159: code <= 5;
				 160: code <= 0;
				 161: code <= 2;
				 162: code <= 8;
				 163: code <= 4;
				 164: code <= 1;
				 165: code <= 0;
				 166: code <= 2;
				 167: code <= 7;
				 168: code <= 0;
				 169: code <= 1;
				 170: code <= 9;
				 171: code <= 3;
				 172: code <= 8;
				 173: code <= 5;
				 174: code <= 2;
				 175: code <= 1;
				 176: code <= 1;
				 177: code <= 0;
				 178: code <= 5;
				 179: code <= 5;
				 180: code <= 5;
				 181: code <= 9;
				 182: code <= 6;
				 183: code <= 4;
				 184: code <= 4;
				 185: code <= 6;
				 186: code <= 2;
				 187: code <= 2;
				 188: code <= 9;
				 189: code <= 4;
				 190: code <= 8;
				 191: code <= 9;
				 192: code <= 5;
				 193: code <= 4;
				 194: code <= 9;
				 195: code <= 3;
				 196: code <= 0;
				 197: code <= 3;
				 198: code <= 8;
				 199: code <= 1;
				 200: code <= 9;
				 201: code <= 6;
				 202: code <= 4;
				 203: code <= 4;
				 204: code <= 2;
				 205: code <= 8;
				 206: code <= 8;
				 207: code <= 1;
				 208: code <= 0;
				 209: code <= 9;
				 210: code <= 7;
				 211: code <= 5;
				 212: code <= 6;
				 213: code <= 6;
				 214: code <= 5;
				 215: code <= 9;
				 216: code <= 3;
				 217: code <= 3;
				 218: code <= 4;
				 219: code <= 4;
				 220: code <= 6;
				 221: code <= 1;
				 222: code <= 2;
				 223: code <= 8;
				 224: code <= 4;
				 225: code <= 7;
				 226: code <= 5;
				 227: code <= 6;
				 228: code <= 4;
				 229: code <= 8;
				 230: code <= 2;
				 231: code <= 3;
				 232: code <= 3;
				 233: code <= 7;
				 234: code <= 8;
				 235: code <= 6;
				 236: code <= 7;
				 237: code <= 8;
				 238: code <= 3;
				 239: code <= 1;
				 240: code <= 6;
				 241: code <= 5;
				 242: code <= 2;
				 243: code <= 7;
				 244: code <= 1;
				 245: code <= 2;
				 246: code <= 0;
				 247: code <= 1;
				 248: code <= 9;
				 249: code <= 0;
				 250: code <= 9;
				 251: code <= 1;
				 252: code <= 4;
				 253: code <= 5;
				 254: code <= 6;
				 255: code <= 4;
				 256: code <= 8;
				 257: code <= 5;
				 258: code <= 6;
				 259: code <= 6;
				 260: code <= 9;
				 261: code <= 2;
				 262: code <= 3;
				 263: code <= 4;
				 264: code <= 6;
				 265: code <= 0;
				 266: code <= 3;
				 267: code <= 4;
				 268: code <= 8;
				 269: code <= 6;
				 270: code <= 1;
				 271: code <= 0;
				 272: code <= 4;
				 273: code <= 5;
				 274: code <= 4;
				 275: code <= 3;
				 276: code <= 2;
				 277: code <= 6;
				 278: code <= 6;
				 279: code <= 4;
				 280: code <= 8;
				 281: code <= 2;
				 282: code <= 1;
				 283: code <= 3;
				 284: code <= 3;
				 285: code <= 9;
				 286: code <= 3;
				 287: code <= 6;
				 288: code <= 0;
				 289: code <= 7;
				 290: code <= 2;
				 291: code <= 6;
				 292: code <= 0;
				 293: code <= 2;
				 294: code <= 4;
				 295: code <= 9;
				 296: code <= 1;
				 297: code <= 4;
				 298: code <= 1;
				 299: code <= 2;
				 300: code <= 7;
				 301: code <= 3;
				 302: code <= 7;
				 303: code <= 2;
				 304: code <= 4;
				 305: code <= 5;
				 306: code <= 8;
				 307: code <= 7;
				 308: code <= 0;
				 309: code <= 0;
				 310: code <= 6;
				 311: code <= 6;
				 312: code <= 0;
				 313: code <= 6;
				 314: code <= 3;
				 315: code <= 1;
				 316: code <= 5;
				 317: code <= 5;
				 318: code <= 8;
				 319: code <= 8;
				 320: code <= 1;
				 321: code <= 7;
				 322: code <= 4;
				 323: code <= 8;
				 324: code <= 8;
				 325: code <= 1;
				 326: code <= 5;
				 327: code <= 2;
				 328: code <= 0;
				 329: code <= 9;
				 330: code <= 2;
				 331: code <= 0;
				 332: code <= 9;
				 333: code <= 6;
				 334: code <= 2;
				 335: code <= 8;
				 336: code <= 2;
				 337: code <= 9;
				 338: code <= 2;
				 339: code <= 5;
				 340: code <= 4;
				 341: code <= 0;
				 342: code <= 9;
				 343: code <= 1;
				 344: code <= 7;
				 345: code <= 1;
				 346: code <= 5;
				 347: code <= 3;
				 348: code <= 6;
				 349: code <= 4;
				 350: code <= 3;
				 351: code <= 6;
				 352: code <= 7;
				 353: code <= 8;
				 354: code <= 9;
				 355: code <= 2;
				 356: code <= 5;
				 357: code <= 9;
				 358: code <= 0;
				 359: code <= 3;
				 360: code <= 6;
				 361: code <= 0;
				 362: code <= 0;
				 363: code <= 1;
				 364: code <= 1;
				 365: code <= 3;
				 366: code <= 3;
				 367: code <= 0;
				 368: code <= 5;
				 369: code <= 3;
				 370: code <= 0;
				 371: code <= 5;
				 372: code <= 4;
				 373: code <= 8;
				 374: code <= 8;
				 375: code <= 2;
				 376: code <= 0;
				 377: code <= 4;
				 378: code <= 6;
				 379: code <= 6;
				 380: code <= 5;
				 381: code <= 2;
				 382: code <= 1;
				 383: code <= 3;
				 384: code <= 8;
				 385: code <= 4;
				 386: code <= 1;
				 387: code <= 4;
				 388: code <= 6;
				 389: code <= 9;
				 390: code <= 5;
				 391: code <= 1;
				 392: code <= 9;
				 393: code <= 4;
				 394: code <= 1;
				 395: code <= 5;
				 396: code <= 1;
				 397: code <= 1;
				 398: code <= 6;
				 399: code <= 0;
				 400: code <= 9;
				 401: code <= 4;
				 402: code <= 3;
				 403: code <= 3;
				 404: code <= 0;
				 405: code <= 5;
				 406: code <= 7;
				 407: code <= 2;
				 408: code <= 7;
				 409: code <= 0;
				 410: code <= 3;
				 411: code <= 6;
				 412: code <= 5;
				 413: code <= 7;
				 414: code <= 5;
				 415: code <= 9;
				 416: code <= 5;
				 417: code <= 9;
				 418: code <= 1;
				 419: code <= 9;
				 420: code <= 5;
				 421: code <= 3;
				 422: code <= 0;
				 423: code <= 9;
				 424: code <= 2;
				 425: code <= 1;
				 426: code <= 8;
				 427: code <= 6;
				 428: code <= 1;
				 429: code <= 1;
				 430: code <= 7;
				 431: code <= 3;
				 432: code <= 8;
				 433: code <= 1;
				 434: code <= 9;
				 435: code <= 3;
				 436: code <= 2;
				 437: code <= 6;
				 438: code <= 1;
				 439: code <= 1;
				 440: code <= 7;
				 441: code <= 9;
				 442: code <= 3;
				 443: code <= 1;
				 444: code <= 0;
				 445: code <= 5;
				 446: code <= 1;
				 447: code <= 1;
				 448: code <= 8;
				 449: code <= 5;
				 450: code <= 4;
				 451: code <= 8;
				 452: code <= 0;
				 453: code <= 7;
				 454: code <= 4;
				 455: code <= 4;
				 456: code <= 6;
				 457: code <= 2;
				 458: code <= 3;
				 459: code <= 7;
				 460: code <= 9;
				 461: code <= 9;
				 462: code <= 6;
				 463: code <= 2;
				 464: code <= 7;
				 465: code <= 4;
				 466: code <= 9;
				 467: code <= 5;
				 468: code <= 6;
				 469: code <= 7;
				 470: code <= 3;
				 471: code <= 5;
				 472: code <= 1;
				 473: code <= 8;
				 474: code <= 8;
				 475: code <= 5;
				 476: code <= 7;
				 477: code <= 5;
				 478: code <= 2;
				 479: code <= 7;
				 480: code <= 2;
				 481: code <= 4;
				 482: code <= 8;
				 483: code <= 9;
				 484: code <= 1;
				 485: code <= 2;
				 486: code <= 2;
				 487: code <= 7;
				 488: code <= 9;
				 489: code <= 3;
				 490: code <= 8;
				 491: code <= 1;
				 492: code <= 8;
				 493: code <= 3;
				 494: code <= 0;
				 495: code <= 1;
				 496: code <= 1;
				 497: code <= 9;
				 498: code <= 4;
				 499: code <= 9;
				 500: code <= 1;
				 501: code <= 2;
				 502: code <= 9;
				 503: code <= 8;
				 504: code <= 3;
				 505: code <= 3;
				 506: code <= 6;
				 507: code <= 7;
				 508: code <= 3;
				 509: code <= 3;
				 510: code <= 6;
				 511: code <= 2;
				 512: code <= 4;
				 513: code <= 4;
				 514: code <= 0;
				 515: code <= 6;
				 516: code <= 5;
				 517: code <= 6;
				 518: code <= 6;
				 519: code <= 4;
				 520: code <= 3;
				 521: code <= 0;
				 522: code <= 8;
				 523: code <= 6;
				 524: code <= 0;
				 525: code <= 2;
				 526: code <= 1;
				 527: code <= 3;
				 528: code <= 9;
				 529: code <= 4;
				 530: code <= 9;
				 531: code <= 4;
				 532: code <= 6;
				 533: code <= 3;
				 534: code <= 9;
				 535: code <= 5;
				 536: code <= 2;
				 537: code <= 2;
				 538: code <= 4;
				 539: code <= 7;
				 540: code <= 3;
				 541: code <= 7;
				 542: code <= 1;
				 543: code <= 9;
				 544: code <= 0;
				 545: code <= 7;
				 546: code <= 0;
				 547: code <= 2;
				 548: code <= 1;
				 549: code <= 7;
				 550: code <= 9;
				 551: code <= 8;
				 552: code <= 6;
				 553: code <= 0;
				 554: code <= 9;
				 555: code <= 4;
				 556: code <= 3;
				 557: code <= 7;
				 558: code <= 0;
				 559: code <= 2;
				 560: code <= 7;
				 561: code <= 7;
				 562: code <= 0;
				 563: code <= 5;
				 564: code <= 3;
				 565: code <= 9;
				 566: code <= 2;
				 567: code <= 1;
				 568: code <= 7;
				 569: code <= 1;
				 570: code <= 7;
				 571: code <= 6;
				 572: code <= 2;
				 573: code <= 9;
				 574: code <= 3;
				 575: code <= 1;
				 576: code <= 7;
				 577: code <= 6;
				 578: code <= 7;
				 579: code <= 5;
				 580: code <= 2;
				 581: code <= 3;
				 582: code <= 8;
				 583: code <= 4;
				 584: code <= 6;
				 585: code <= 7;
				 586: code <= 4;
				 587: code <= 8;
				 588: code <= 1;
				 589: code <= 8;
				 590: code <= 4;
				 591: code <= 6;
				 592: code <= 7;
				 593: code <= 6;
				 594: code <= 6;
				 595: code <= 9;
				 596: code <= 4;
				 597: code <= 0;
				 598: code <= 5;
				 599: code <= 1;
				 600: code <= 3;
				 601: code <= 2;
				 602: code <= 0;
				 603: code <= 0;
				 604: code <= 0;
				 605: code <= 5;
				 606: code <= 6;
				 607: code <= 8;
				 608: code <= 1;
				 609: code <= 2;
				 610: code <= 7;
				 611: code <= 1;
				 612: code <= 4;
				 613: code <= 5;
				 614: code <= 2;
				 615: code <= 6;
				 616: code <= 3;
				 617: code <= 5;
				 618: code <= 6;
				 619: code <= 0;
				 620: code <= 8;
				 621: code <= 2;
				 622: code <= 7;
				 623: code <= 7;
				 624: code <= 8;
				 625: code <= 5;
				 626: code <= 7;
				 627: code <= 7;
				 628: code <= 1;
				 629: code <= 3;
				 630: code <= 4;
				 631: code <= 2;
				 632: code <= 7;
				 633: code <= 5;
				 634: code <= 7;
				 635: code <= 7;
				 636: code <= 8;
				 637: code <= 9;
				 638: code <= 6;
				 639: code <= 0;
				 640: code <= 9;
				 641: code <= 1;
				 642: code <= 7;
				 643: code <= 3;
				 644: code <= 6;
				 645: code <= 3;
				 646: code <= 7;
				 647: code <= 1;
				 648: code <= 7;
				 649: code <= 8;
				 650: code <= 7;
				 651: code <= 2;
				 652: code <= 1;
				 653: code <= 4;
				 654: code <= 6;
				 655: code <= 8;
				 656: code <= 4;
				 657: code <= 4;
				 658: code <= 0;
				 659: code <= 9;
				 660: code <= 0;
				 661: code <= 1;
				 662: code <= 2;
				 663: code <= 2;
				 664: code <= 4;
				 665: code <= 9;
				 666: code <= 5;
				 667: code <= 3;
				 668: code <= 4;
				 669: code <= 3;
				 670: code <= 0;
				 671: code <= 1;
				 672: code <= 4;
				 673: code <= 6;
				 674: code <= 5;
				 675: code <= 4;
				 676: code <= 9;
				 677: code <= 5;
				 678: code <= 8;
				 679: code <= 5;
				 680: code <= 3;
				 681: code <= 7;
				 682: code <= 1;
				 683: code <= 0;
				 684: code <= 5;
				 685: code <= 0;
				 686: code <= 7;
				 687: code <= 9;
				 688: code <= 2;
				 689: code <= 2;
				 690: code <= 7;
				 691: code <= 9;
				 692: code <= 6;
				 693: code <= 8;
				 694: code <= 9;
				 695: code <= 2;
				 696: code <= 5;
				 697: code <= 8;
				 698: code <= 9;
				 699: code <= 2;
				 700: code <= 3;
				 701: code <= 5;
				 702: code <= 4;
				 703: code <= 2;
				 704: code <= 0;
				 705: code <= 1;
				 706: code <= 9;
				 707: code <= 9;
				 708: code <= 5;
				 709: code <= 6;
				 710: code <= 1;
				 711: code <= 1;
				 712: code <= 2;
				 713: code <= 1;
				 714: code <= 2;
				 715: code <= 9;
				 716: code <= 0;
				 717: code <= 2;
				 718: code <= 1;
				 719: code <= 9;
				 720: code <= 6;
				 721: code <= 0;
				 722: code <= 8;
				 723: code <= 6;
				 724: code <= 4;
				 725: code <= 0;
				 726: code <= 3;
				 727: code <= 4;
				 728: code <= 4;
				 729: code <= 1;
				 730: code <= 8;
				 731: code <= 1;
				 732: code <= 5;
				 733: code <= 9;
				 734: code <= 8;
				 735: code <= 1;
				 736: code <= 3;
				 737: code <= 6;
				 738: code <= 2;
				 739: code <= 9;
				 740: code <= 7;
				 741: code <= 7;
				 742: code <= 4;
				 743: code <= 7;
				 744: code <= 7;
				 745: code <= 1;
				 746: code <= 3;
				 747: code <= 0;
				 748: code <= 9;
				 749: code <= 9;
				 750: code <= 6;
				 751: code <= 0;
				 752: code <= 5;
				 753: code <= 1;
				 754: code <= 8;
				 755: code <= 7;
				 756: code <= 0;
				 757: code <= 7;
				 758: code <= 2;
				 759: code <= 1;
				 760: code <= 1;
				 761: code <= 3;
				 762: code <= 4;
				 763: code <= 9;
				 764: code <= 9;
				 765: code <= 9;
				 766: code <= 9;
				 767: code <= 9;
				 768: code <= 9;
				 769: code <= 8;
				 770: code <= 3;
				 771: code <= 7;
				 772: code <= 2;
				 773: code <= 9;
				 774: code <= 7;
				 775: code <= 8;
				 776: code <= 0;
				 777: code <= 4;
				 778: code <= 9;
				 779: code <= 9;
				 780: code <= 5;
				 781: code <= 1;
				 782: code <= 0;
				 783: code <= 5;
				 784: code <= 9;
				 785: code <= 7;
				 786: code <= 3;
				 787: code <= 1;
				 788: code <= 7;
				 789: code <= 3;
				 790: code <= 2;
				 791: code <= 8;
				 792: code <= 1;
				 793: code <= 6;
				 794: code <= 0;
				 795: code <= 9;
				 796: code <= 6;
				 797: code <= 3;
				 798: code <= 1;
				 799: code <= 8;
				 800: code <= 5;
				 801: code <= 9;
				 802: code <= 5;
				 803: code <= 0;
				 804: code <= 2;
				 805: code <= 4;
				 806: code <= 4;
				 807: code <= 5;
				 808: code <= 9;
				 809: code <= 4;
				 810: code <= 5;
				 811: code <= 5;
				 812: code <= 3;
				 813: code <= 4;
				 814: code <= 6;
				 815: code <= 9;
				 816: code <= 0;
				 817: code <= 8;
				 818: code <= 3;
				 819: code <= 0;
				 820: code <= 2;
				 821: code <= 6;
				 822: code <= 4;
				 823: code <= 2;
				 824: code <= 5;
				 825: code <= 2;
				 826: code <= 2;
				 827: code <= 3;
				 828: code <= 0;
				 829: code <= 8;
				 830: code <= 2;
				 831: code <= 5;
				 832: code <= 3;
				 833: code <= 3;
				 834: code <= 4;
				 835: code <= 4;
				 836: code <= 6;
				 837: code <= 8;
				 838: code <= 5;
				 839: code <= 0;
				 840: code <= 3;
				 841: code <= 5;
				 842: code <= 2;
				 843: code <= 6;
				 844: code <= 1;
				 845: code <= 9;
				 846: code <= 3;
				 847: code <= 1;
				 848: code <= 1;
				 849: code <= 8;
				 850: code <= 8;
				 851: code <= 1;
				 852: code <= 7;
				 853: code <= 1;
				 854: code <= 0;
				 855: code <= 1;
				 856: code <= 0;
				 857: code <= 0;
				 858: code <= 0;
				 859: code <= 3;
				 860: code <= 1;
				 861: code <= 3;
				 862: code <= 7;
				 863: code <= 8;
				 864: code <= 3;
				 865: code <= 8;
				 866: code <= 7;
				 867: code <= 5;
				 868: code <= 2;
				 869: code <= 8;
				 870: code <= 8;
				 871: code <= 6;
				 872: code <= 5;
				 873: code <= 8;
				 874: code <= 7;
				 875: code <= 5;
				 876: code <= 3;
				 877: code <= 3;
				 878: code <= 2;
				 879: code <= 0;
				 880: code <= 8;
				 881: code <= 3;
				 882: code <= 8;
				 883: code <= 1;
				 884: code <= 4;
				 885: code <= 2;
				 886: code <= 0;
				 887: code <= 6;
				 888: code <= 1;
				 889: code <= 7;
				 890: code <= 1;
				 891: code <= 7;
				 892: code <= 7;
				 893: code <= 6;
				 894: code <= 6;
				 895: code <= 9;
				 896: code <= 1;
				 897: code <= 4;
				 898: code <= 7;
				 899: code <= 3;
				 900: code <= 0;
				 901: code <= 3;
				 902: code <= 5;
				 903: code <= 9;
				 904: code <= 8;
				 905: code <= 2;
				 906: code <= 5;
				 907: code <= 3;
				 908: code <= 4;
				 909: code <= 9;
				 910: code <= 0;
				 911: code <= 4;
				 912: code <= 2;
				 913: code <= 8;
				 914: code <= 7;
				 915: code <= 5;
				 916: code <= 5;
				 917: code <= 4;
				 918: code <= 6;
				 919: code <= 8;
				 920: code <= 7;
				 921: code <= 3;
				 922: code <= 1;
				 923: code <= 1;
				 924: code <= 5;
				 925: code <= 9;
				 926: code <= 5;
				 927: code <= 6;
				 928: code <= 2;
				 929: code <= 8;
				 930: code <= 6;
				 931: code <= 3;
				 932: code <= 8;
				 933: code <= 8;
				 934: code <= 2;
				 935: code <= 3;
				 936: code <= 5;
				 937: code <= 3;
				 938: code <= 7;
				 939: code <= 8;
				 940: code <= 7;
				 941: code <= 5;
				 942: code <= 9;
				 943: code <= 3;
				 944: code <= 7;
				 945: code <= 5;
				 946: code <= 1;
				 947: code <= 9;
				 948: code <= 5;
				 949: code <= 7;
				 950: code <= 7;
				 951: code <= 8;
				 952: code <= 1;
				 953: code <= 8;
				 954: code <= 5;
				 955: code <= 7;
				 956: code <= 7;
				 957: code <= 8;
				 958: code <= 0;
				 959: code <= 5;
				 960: code <= 3;
				 961: code <= 2;
				 962: code <= 1;
				 963: code <= 7;
				 964: code <= 1;
				 965: code <= 2;
				 966: code <= 2;
				 967: code <= 6;
				 968: code <= 8;
				 969: code <= 0;
				 970: code <= 6;
				 971: code <= 6;
				 972: code <= 1;
				 973: code <= 3;
				 974: code <= 0;
				 975: code <= 0;
				 976: code <= 1;
				 977: code <= 9;
				 978: code <= 2;
				 979: code <= 7;
				 980: code <= 8;
				 981: code <= 7;
				 982: code <= 6;
				 983: code <= 6;
				 984: code <= 1;
				 985: code <= 1;
				 986: code <= 1;
				 987: code <= 9;
				 988: code <= 5;
				 989: code <= 9;
				 990: code <= 0;
				 991: code <= 9;
				 992: code <= 2;
				 993: code <= 1;
				 994: code <= 6;
				 995: code <= 4;
				 996: code <= 2;
				 997: code <= 0;
				 998: code <= 1;
				 999: code <= 9;
				1000: code <= 8;
				1001: code <= 9;
				1002: code <= 3;
				1003: code <= 8;
				1004: code <= 0;
				1005: code <= 9;
				1006: code <= 5;
				1007: code <= 2;
				1008: code <= 5;
				1009: code <= 7;
				1010: code <= 2;
				1011: code <= 0;
				1012: code <= 1;
				1013: code <= 0;
				1014: code <= 6;
				1015: code <= 5;
				1016: code <= 4;
				1017: code <= 8;
				1018: code <= 5;
				1019: code <= 8;
				1020: code <= 6;
				1021: code <= 3;
				1022: code <= 2;
				1023: code <= 7;
			endcase
		end
	end

	decoder decoder(.code(code), .segments(led_out));

endmodule

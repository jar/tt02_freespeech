module jar_pi
(
	input  [7:0] io_in,
	output [7:0] io_out
);
	wire       clk      = io_in[0];
	wire       reset    = io_in[1];
	//wire       stream   = io_in[2];
	wire [4:0] io_index = io_in[7:3];

	reg [9:0] index;
	reg [3:0] code;

	always @(posedge clk) begin
		if (reset) begin
			index <= {io_index, index[9:5]};
		end
		else begin //if (stream) begin
			index <= index + 1;

			/* verilator lint_off CASEX */
			casex(index)
				0: code <= 4'bx011;
				1: code <= 4'b1010;
				2: code <= 4'b0001;
				3: code <= 4'bx100;
				4: code <= 4'b0001;
				5: code <= 4'bx101;
				6: code <= 4'b1001;
				7: code <= 4'b0010;
				8: code <= 4'bx110;
				9: code <= 4'bx101;
				10: code <= 4'bx011;
				11: code <= 4'bx101;
				12: code <= 4'b1000;
				13: code <= 4'b1001;
				14: code <= 4'bx111;
				15: code <= 4'b1001;
				16: code <= 4'bx011;
				17: code <= 4'b0010;
				18: code <= 4'bx011;
				19: code <= 4'b1000;
				20: code <= 4'bx100;
				21: code <= 4'bx110;
				22: code <= 4'b0010;
				23: code <= 4'bx110;
				24: code <= 4'bx100;
				25: code <= 4'bx011;
				26: code <= 4'bx011;
				27: code <= 4'b1000;
				28: code <= 4'bx011;
				29: code <= 4'b0010;
				30: code <= 4'bx111;
				31: code <= 4'b1001;
				32: code <= 4'bx101;
				33: code <= 4'b0000;
				34: code <= 4'b0010;
				35: code <= 4'b1000;
				36: code <= 4'b1000;
				37: code <= 4'bx100;
				38: code <= 4'b0001;
				39: code <= 4'b1001;
				40: code <= 4'bx111;
				41: code <= 4'b0001;
				42: code <= 4'bx110;
				43: code <= 4'b1001;
				44: code <= 4'bx011;
				45: code <= 4'b1001;
				46: code <= 4'b1001;
				47: code <= 4'bx011;
				48: code <= 4'bx111;
				49: code <= 4'bx101;
				50: code <= 4'b0001;
				51: code <= 4'b0000;
				52: code <= 4'bx101;
				53: code <= 4'b1000;
				54: code <= 4'b0010;
				55: code <= 4'b0000;
				56: code <= 4'b1001;
				57: code <= 4'bx111;
				58: code <= 4'bx100;
				59: code <= 4'b1001;
				60: code <= 4'bx100;
				61: code <= 4'bx100;
				62: code <= 4'bx101;
				63: code <= 4'b1001;
				64: code <= 4'b0010;
				65: code <= 4'bx011;
				66: code <= 4'b0000;
				67: code <= 4'bx111;
				68: code <= 4'b1000;
				69: code <= 4'b0001;
				70: code <= 4'bx110;
				71: code <= 4'bx100;
				72: code <= 4'b0000;
				73: code <= 4'bx110;
				74: code <= 4'b0010;
				75: code <= 4'b1000;
				76: code <= 4'bx110;
				77: code <= 4'b0010;
				78: code <= 4'b0000;
				79: code <= 4'b1000;
				80: code <= 4'b1001;
				81: code <= 4'b1001;
				82: code <= 4'b1000;
				83: code <= 4'bx110;
				84: code <= 4'b0010;
				85: code <= 4'b1000;
				86: code <= 4'b0000;
				87: code <= 4'bx011;
				88: code <= 4'bx100;
				89: code <= 4'b1000;
				90: code <= 4'b0010;
				91: code <= 4'bx101;
				92: code <= 4'bx011;
				93: code <= 4'bx100;
				94: code <= 4'b0010;
				95: code <= 4'b0001;
				96: code <= 4'b0001;
				97: code <= 4'bx111;
				98: code <= 4'b0000;
				99: code <= 4'bx110;
				100: code <= 4'bx111;
				101: code <= 4'b1001;
				102: code <= 4'b1000;
				103: code <= 4'b0010;
				104: code <= 4'b0001;
				105: code <= 4'bx100;
				106: code <= 4'b1000;
				107: code <= 4'b0000;
				108: code <= 4'b1000;
				109: code <= 4'bx110;
				110: code <= 4'bx101;
				111: code <= 4'b0001;
				112: code <= 4'bx011;
				113: code <= 4'b0010;
				114: code <= 4'b1000;
				115: code <= 4'b0010;
				116: code <= 4'bx011;
				117: code <= 4'b0000;
				118: code <= 4'bx110;
				119: code <= 4'bx110;
				120: code <= 4'bx100;
				121: code <= 4'bx111;
				122: code <= 4'b0000;
				123: code <= 4'b1001;
				124: code <= 4'bx011;
				125: code <= 4'b1000;
				126: code <= 4'bx100;
				127: code <= 4'bx100;
				128: code <= 4'bx110;
				129: code <= 4'b0000;
				130: code <= 4'b1001;
				131: code <= 4'bx101;
				132: code <= 4'bx101;
				133: code <= 4'b0000;
				134: code <= 4'bx101;
				135: code <= 4'b1000;
				136: code <= 4'b0010;
				137: code <= 4'b0010;
				138: code <= 4'bx011;
				139: code <= 4'b0001;
				140: code <= 4'bx111;
				141: code <= 4'b0010;
				142: code <= 4'bx101;
				143: code <= 4'bx011;
				144: code <= 4'bx101;
				145: code <= 4'b1001;
				146: code <= 4'bx100;
				147: code <= 4'b0000;
				148: code <= 4'b1000;
				149: code <= 4'b0001;
				150: code <= 4'b0010;
				151: code <= 4'b1000;
				152: code <= 4'bx100;
				153: code <= 4'b1000;
				154: code <= 4'b0001;
				155: code <= 4'b0001;
				156: code <= 4'b0001;
				157: code <= 4'bx111;
				158: code <= 4'bx100;
				159: code <= 4'bx101;
				160: code <= 4'b0000;
				161: code <= 4'b0010;
				162: code <= 4'b1000;
				163: code <= 4'bx100;
				164: code <= 4'b0001;
				165: code <= 4'b0000;
				166: code <= 4'b0010;
				167: code <= 4'bx111;
				168: code <= 4'b0000;
				169: code <= 4'b0001;
				170: code <= 4'b1001;
				171: code <= 4'bx011;
				172: code <= 4'b1000;
				173: code <= 4'bx101;
				174: code <= 4'b0010;
				175: code <= 4'b0001;
				176: code <= 4'b0001;
				177: code <= 4'b0000;
				178: code <= 4'bx101;
				179: code <= 4'bx101;
				180: code <= 4'bx101;
				181: code <= 4'b1001;
				182: code <= 4'bx110;
				183: code <= 4'bx100;
				184: code <= 4'bx100;
				185: code <= 4'bx110;
				186: code <= 4'b0010;
				187: code <= 4'b0010;
				188: code <= 4'b1001;
				189: code <= 4'bx100;
				190: code <= 4'b1000;
				191: code <= 4'b1001;
				192: code <= 4'bx101;
				193: code <= 4'bx100;
				194: code <= 4'b1001;
				195: code <= 4'bx011;
				196: code <= 4'b0000;
				197: code <= 4'bx011;
				198: code <= 4'b1000;
				199: code <= 4'b0001;
				200: code <= 4'b1001;
				201: code <= 4'bx110;
				202: code <= 4'bx100;
				203: code <= 4'bx100;
				204: code <= 4'b0010;
				205: code <= 4'b1000;
				206: code <= 4'b1000;
				207: code <= 4'b0001;
				208: code <= 4'b0000;
				209: code <= 4'b1001;
				210: code <= 4'bx111;
				211: code <= 4'bx101;
				212: code <= 4'bx110;
				213: code <= 4'bx110;
				214: code <= 4'bx101;
				215: code <= 4'b1001;
				216: code <= 4'bx011;
				217: code <= 4'bx011;
				218: code <= 4'bx100;
				219: code <= 4'bx100;
				220: code <= 4'bx110;
				221: code <= 4'b0001;
				222: code <= 4'b0010;
				223: code <= 4'b1000;
				224: code <= 4'bx100;
				225: code <= 4'bx111;
				226: code <= 4'bx101;
				227: code <= 4'bx110;
				228: code <= 4'bx100;
				229: code <= 4'b1000;
				230: code <= 4'b0010;
				231: code <= 4'bx011;
				232: code <= 4'bx011;
				233: code <= 4'bx111;
				234: code <= 4'b1000;
				235: code <= 4'bx110;
				236: code <= 4'bx111;
				237: code <= 4'b1000;
				238: code <= 4'bx011;
				239: code <= 4'b0001;
				240: code <= 4'bx110;
				241: code <= 4'bx101;
				242: code <= 4'b0010;
				243: code <= 4'bx111;
				244: code <= 4'b0001;
				245: code <= 4'b0010;
				246: code <= 4'b0000;
				247: code <= 4'b0001;
				248: code <= 4'b1001;
				249: code <= 4'b0000;
				250: code <= 4'b1001;
				251: code <= 4'b0001;
				252: code <= 4'bx100;
				253: code <= 4'bx101;
				254: code <= 4'bx110;
				255: code <= 4'bx100;
				256: code <= 4'b1000;
				257: code <= 4'bx101;
				258: code <= 4'bx110;
				259: code <= 4'bx110;
				260: code <= 4'b1001;
				261: code <= 4'b0010;
				262: code <= 4'bx011;
				263: code <= 4'bx100;
				264: code <= 4'bx110;
				265: code <= 4'b0000;
				266: code <= 4'bx011;
				267: code <= 4'bx100;
				268: code <= 4'b1000;
				269: code <= 4'bx110;
				270: code <= 4'b0001;
				271: code <= 4'b0000;
				272: code <= 4'bx100;
				273: code <= 4'bx101;
				274: code <= 4'bx100;
				275: code <= 4'bx011;
				276: code <= 4'b0010;
				277: code <= 4'bx110;
				278: code <= 4'bx110;
				279: code <= 4'bx100;
				280: code <= 4'b1000;
				281: code <= 4'b0010;
				282: code <= 4'b0001;
				283: code <= 4'bx011;
				284: code <= 4'bx011;
				285: code <= 4'b1001;
				286: code <= 4'bx011;
				287: code <= 4'bx110;
				288: code <= 4'b0000;
				289: code <= 4'bx111;
				290: code <= 4'b0010;
				291: code <= 4'bx110;
				292: code <= 4'b0000;
				293: code <= 4'b0010;
				294: code <= 4'bx100;
				295: code <= 4'b1001;
				296: code <= 4'b0001;
				297: code <= 4'bx100;
				298: code <= 4'b0001;
				299: code <= 4'b0010;
				300: code <= 4'bx111;
				301: code <= 4'bx011;
				302: code <= 4'bx111;
				303: code <= 4'b0010;
				304: code <= 4'bx100;
				305: code <= 4'bx101;
				306: code <= 4'b1000;
				307: code <= 4'bx111;
				308: code <= 4'b0000;
				309: code <= 4'b0000;
				310: code <= 4'bx110;
				311: code <= 4'bx110;
				312: code <= 4'b0000;
				313: code <= 4'bx110;
				314: code <= 4'bx011;
				315: code <= 4'b0001;
				316: code <= 4'bx101;
				317: code <= 4'bx101;
				318: code <= 4'b1000;
				319: code <= 4'b1000;
				320: code <= 4'b0001;
				321: code <= 4'bx111;
				322: code <= 4'bx100;
				323: code <= 4'b1000;
				324: code <= 4'b1000;
				325: code <= 4'b0001;
				326: code <= 4'bx101;
				327: code <= 4'b0010;
				328: code <= 4'b0000;
				329: code <= 4'b1001;
				330: code <= 4'b0010;
				331: code <= 4'b0000;
				332: code <= 4'b1001;
				333: code <= 4'bx110;
				334: code <= 4'b0010;
				335: code <= 4'b1000;
				336: code <= 4'b0010;
				337: code <= 4'b1001;
				338: code <= 4'b0010;
				339: code <= 4'bx101;
				340: code <= 4'bx100;
				341: code <= 4'b0000;
				342: code <= 4'b1001;
				343: code <= 4'b0001;
				344: code <= 4'bx111;
				345: code <= 4'b0001;
				346: code <= 4'bx101;
				347: code <= 4'bx011;
				348: code <= 4'bx110;
				349: code <= 4'bx100;
				350: code <= 4'bx011;
				351: code <= 4'bx110;
				352: code <= 4'bx111;
				353: code <= 4'b1000;
				354: code <= 4'b1001;
				355: code <= 4'b0010;
				356: code <= 4'bx101;
				357: code <= 4'b1001;
				358: code <= 4'b0000;
				359: code <= 4'bx011;
				360: code <= 4'bx110;
				361: code <= 4'b0000;
				362: code <= 4'b0000;
				363: code <= 4'b0001;
				364: code <= 4'b0001;
				365: code <= 4'bx011;
				366: code <= 4'bx011;
				367: code <= 4'b0000;
				368: code <= 4'bx101;
				369: code <= 4'bx011;
				370: code <= 4'b0000;
				371: code <= 4'bx101;
				372: code <= 4'bx100;
				373: code <= 4'b1000;
				374: code <= 4'b1000;
				375: code <= 4'b0010;
				376: code <= 4'b0000;
				377: code <= 4'bx100;
				378: code <= 4'bx110;
				379: code <= 4'bx110;
				380: code <= 4'bx101;
				381: code <= 4'b0010;
				382: code <= 4'b0001;
				383: code <= 4'bx011;
				384: code <= 4'b1000;
				385: code <= 4'bx100;
				386: code <= 4'b0001;
				387: code <= 4'bx100;
				388: code <= 4'bx110;
				389: code <= 4'b1001;
				390: code <= 4'bx101;
				391: code <= 4'b0001;
				392: code <= 4'b1001;
				393: code <= 4'bx100;
				394: code <= 4'b0001;
				395: code <= 4'bx101;
				396: code <= 4'b0001;
				397: code <= 4'b0001;
				398: code <= 4'bx110;
				399: code <= 4'b0000;
				400: code <= 4'b1001;
				401: code <= 4'bx100;
				402: code <= 4'bx011;
				403: code <= 4'bx011;
				404: code <= 4'b0000;
				405: code <= 4'bx101;
				406: code <= 4'bx111;
				407: code <= 4'b0010;
				408: code <= 4'bx111;
				409: code <= 4'b0000;
				410: code <= 4'bx011;
				411: code <= 4'bx110;
				412: code <= 4'bx101;
				413: code <= 4'bx111;
				414: code <= 4'bx101;
				415: code <= 4'b1001;
				416: code <= 4'bx101;
				417: code <= 4'b1001;
				418: code <= 4'b0001;
				419: code <= 4'b1001;
				420: code <= 4'bx101;
				421: code <= 4'bx011;
				422: code <= 4'b0000;
				423: code <= 4'b1001;
				424: code <= 4'b0010;
				425: code <= 4'b0001;
				426: code <= 4'b1000;
				427: code <= 4'bx110;
				428: code <= 4'b0001;
				429: code <= 4'b0001;
				430: code <= 4'bx111;
				431: code <= 4'bx011;
				432: code <= 4'b1000;
				433: code <= 4'b0001;
				434: code <= 4'b1001;
				435: code <= 4'bx011;
				436: code <= 4'b0010;
				437: code <= 4'bx110;
				438: code <= 4'b0001;
				439: code <= 4'b0001;
				440: code <= 4'bx111;
				441: code <= 4'b1001;
				442: code <= 4'bx011;
				443: code <= 4'b0001;
				444: code <= 4'b0000;
				445: code <= 4'bx101;
				446: code <= 4'b0001;
				447: code <= 4'b0001;
				448: code <= 4'b1000;
				449: code <= 4'bx101;
				450: code <= 4'bx100;
				451: code <= 4'b1000;
				452: code <= 4'b0000;
				453: code <= 4'bx111;
				454: code <= 4'bx100;
				455: code <= 4'bx100;
				456: code <= 4'bx110;
				457: code <= 4'b0010;
				458: code <= 4'bx011;
				459: code <= 4'bx111;
				460: code <= 4'b1001;
				461: code <= 4'b1001;
				462: code <= 4'bx110;
				463: code <= 4'b0010;
				464: code <= 4'bx111;
				465: code <= 4'bx100;
				466: code <= 4'b1001;
				467: code <= 4'bx101;
				468: code <= 4'bx110;
				469: code <= 4'bx111;
				470: code <= 4'bx011;
				471: code <= 4'bx101;
				472: code <= 4'b0001;
				473: code <= 4'b1000;
				474: code <= 4'b1000;
				475: code <= 4'bx101;
				476: code <= 4'bx111;
				477: code <= 4'bx101;
				478: code <= 4'b0010;
				479: code <= 4'bx111;
				480: code <= 4'b0010;
				481: code <= 4'bx100;
				482: code <= 4'b1000;
				483: code <= 4'b1001;
				484: code <= 4'b0001;
				485: code <= 4'b0010;
				486: code <= 4'b0010;
				487: code <= 4'bx111;
				488: code <= 4'b1001;
				489: code <= 4'bx011;
				490: code <= 4'b1000;
				491: code <= 4'b0001;
				492: code <= 4'b1000;
				493: code <= 4'bx011;
				494: code <= 4'b0000;
				495: code <= 4'b0001;
				496: code <= 4'b0001;
				497: code <= 4'b1001;
				498: code <= 4'bx100;
				499: code <= 4'b1001;
				500: code <= 4'b0001;
				501: code <= 4'b0010;
				502: code <= 4'b1001;
				503: code <= 4'b1000;
				504: code <= 4'bx011;
				505: code <= 4'bx011;
				506: code <= 4'bx110;
				507: code <= 4'bx111;
				508: code <= 4'bx011;
				509: code <= 4'bx011;
				510: code <= 4'bx110;
				511: code <= 4'b0010;
				512: code <= 4'bx100;
				513: code <= 4'bx100;
				514: code <= 4'b0000;
				515: code <= 4'bx110;
				516: code <= 4'bx101;
				517: code <= 4'bx110;
				518: code <= 4'bx110;
				519: code <= 4'bx100;
				520: code <= 4'bx011;
				521: code <= 4'b0000;
				522: code <= 4'b1000;
				523: code <= 4'bx110;
				524: code <= 4'b0000;
				525: code <= 4'b0010;
				526: code <= 4'b0001;
				527: code <= 4'bx011;
				528: code <= 4'b1001;
				529: code <= 4'bx100;
				530: code <= 4'b1001;
				531: code <= 4'bx100;
				532: code <= 4'bx110;
				533: code <= 4'bx011;
				534: code <= 4'b1001;
				535: code <= 4'bx101;
				536: code <= 4'b0010;
				537: code <= 4'b0010;
				538: code <= 4'bx100;
				539: code <= 4'bx111;
				540: code <= 4'bx011;
				541: code <= 4'bx111;
				542: code <= 4'b0001;
				543: code <= 4'b1001;
				544: code <= 4'b0000;
				545: code <= 4'bx111;
				546: code <= 4'b0000;
				547: code <= 4'b0010;
				548: code <= 4'b0001;
				549: code <= 4'bx111;
				550: code <= 4'b1001;
				551: code <= 4'b1000;
				552: code <= 4'bx110;
				553: code <= 4'b0000;
				554: code <= 4'b1001;
				555: code <= 4'bx100;
				556: code <= 4'bx011;
				557: code <= 4'bx111;
				558: code <= 4'b0000;
				559: code <= 4'b0010;
				560: code <= 4'bx111;
				561: code <= 4'bx111;
				562: code <= 4'b0000;
				563: code <= 4'bx101;
				564: code <= 4'bx011;
				565: code <= 4'b1001;
				566: code <= 4'b0010;
				567: code <= 4'b0001;
				568: code <= 4'bx111;
				569: code <= 4'b0001;
				570: code <= 4'bx111;
				571: code <= 4'bx110;
				572: code <= 4'b0010;
				573: code <= 4'b1001;
				574: code <= 4'bx011;
				575: code <= 4'b0001;
				576: code <= 4'bx111;
				577: code <= 4'bx110;
				578: code <= 4'bx111;
				579: code <= 4'bx101;
				580: code <= 4'b0010;
				581: code <= 4'bx011;
				582: code <= 4'b1000;
				583: code <= 4'bx100;
				584: code <= 4'bx110;
				585: code <= 4'bx111;
				586: code <= 4'bx100;
				587: code <= 4'b1000;
				588: code <= 4'b0001;
				589: code <= 4'b1000;
				590: code <= 4'bx100;
				591: code <= 4'bx110;
				592: code <= 4'bx111;
				593: code <= 4'bx110;
				594: code <= 4'bx110;
				595: code <= 4'b1001;
				596: code <= 4'bx100;
				597: code <= 4'b0000;
				598: code <= 4'bx101;
				599: code <= 4'b0001;
				600: code <= 4'bx011;
				601: code <= 4'b0010;
				602: code <= 4'b0000;
				603: code <= 4'b0000;
				604: code <= 4'b0000;
				605: code <= 4'bx101;
				606: code <= 4'bx110;
				607: code <= 4'b1000;
				608: code <= 4'b0001;
				609: code <= 4'b0010;
				610: code <= 4'bx111;
				611: code <= 4'b0001;
				612: code <= 4'bx100;
				613: code <= 4'bx101;
				614: code <= 4'b0010;
				615: code <= 4'bx110;
				616: code <= 4'bx011;
				617: code <= 4'bx101;
				618: code <= 4'bx110;
				619: code <= 4'b0000;
				620: code <= 4'b1000;
				621: code <= 4'b0010;
				622: code <= 4'bx111;
				623: code <= 4'bx111;
				624: code <= 4'b1000;
				625: code <= 4'bx101;
				626: code <= 4'bx111;
				627: code <= 4'bx111;
				628: code <= 4'b0001;
				629: code <= 4'bx011;
				630: code <= 4'bx100;
				631: code <= 4'b0010;
				632: code <= 4'bx111;
				633: code <= 4'bx101;
				634: code <= 4'bx111;
				635: code <= 4'bx111;
				636: code <= 4'b1000;
				637: code <= 4'b1001;
				638: code <= 4'bx110;
				639: code <= 4'b0000;
				640: code <= 4'b1001;
				641: code <= 4'b0001;
				642: code <= 4'bx111;
				643: code <= 4'bx011;
				644: code <= 4'bx110;
				645: code <= 4'bx011;
				646: code <= 4'bx111;
				647: code <= 4'b0001;
				648: code <= 4'bx111;
				649: code <= 4'b1000;
				650: code <= 4'bx111;
				651: code <= 4'b0010;
				652: code <= 4'b0001;
				653: code <= 4'bx100;
				654: code <= 4'bx110;
				655: code <= 4'b1000;
				656: code <= 4'bx100;
				657: code <= 4'bx100;
				658: code <= 4'b0000;
				659: code <= 4'b1001;
				660: code <= 4'b0000;
				661: code <= 4'b0001;
				662: code <= 4'b0010;
				663: code <= 4'b0010;
				664: code <= 4'bx100;
				665: code <= 4'b1001;
				666: code <= 4'bx101;
				667: code <= 4'bx011;
				668: code <= 4'bx100;
				669: code <= 4'bx011;
				670: code <= 4'b0000;
				671: code <= 4'b0001;
				672: code <= 4'bx100;
				673: code <= 4'bx110;
				674: code <= 4'bx101;
				675: code <= 4'bx100;
				676: code <= 4'b1001;
				677: code <= 4'bx101;
				678: code <= 4'b1000;
				679: code <= 4'bx101;
				680: code <= 4'bx011;
				681: code <= 4'bx111;
				682: code <= 4'b0001;
				683: code <= 4'b0000;
				684: code <= 4'bx101;
				685: code <= 4'b0000;
				686: code <= 4'bx111;
				687: code <= 4'b1001;
				688: code <= 4'b0010;
				689: code <= 4'b0010;
				690: code <= 4'bx111;
				691: code <= 4'b1001;
				692: code <= 4'bx110;
				693: code <= 4'b1000;
				694: code <= 4'b1001;
				695: code <= 4'b0010;
				696: code <= 4'bx101;
				697: code <= 4'b1000;
				698: code <= 4'b1001;
				699: code <= 4'b0010;
				700: code <= 4'bx011;
				701: code <= 4'bx101;
				702: code <= 4'bx100;
				703: code <= 4'b0010;
				704: code <= 4'b0000;
				705: code <= 4'b0001;
				706: code <= 4'b1001;
				707: code <= 4'b1001;
				708: code <= 4'bx101;
				709: code <= 4'bx110;
				710: code <= 4'b0001;
				711: code <= 4'b0001;
				712: code <= 4'b0010;
				713: code <= 4'b0001;
				714: code <= 4'b0010;
				715: code <= 4'b1001;
				716: code <= 4'b0000;
				717: code <= 4'b0010;
				718: code <= 4'b0001;
				719: code <= 4'b1001;
				720: code <= 4'bx110;
				721: code <= 4'b0000;
				722: code <= 4'b1000;
				723: code <= 4'bx110;
				724: code <= 4'bx100;
				725: code <= 4'b0000;
				726: code <= 4'bx011;
				727: code <= 4'bx100;
				728: code <= 4'bx100;
				729: code <= 4'b0001;
				730: code <= 4'b1000;
				731: code <= 4'b0001;
				732: code <= 4'bx101;
				733: code <= 4'b1001;
				734: code <= 4'b1000;
				735: code <= 4'b0001;
				736: code <= 4'bx011;
				737: code <= 4'bx110;
				738: code <= 4'b0010;
				739: code <= 4'b1001;
				740: code <= 4'bx111;
				741: code <= 4'bx111;
				742: code <= 4'bx100;
				743: code <= 4'bx111;
				744: code <= 4'bx111;
				745: code <= 4'b0001;
				746: code <= 4'bx011;
				747: code <= 4'b0000;
				748: code <= 4'b1001;
				749: code <= 4'b1001;
				750: code <= 4'bx110;
				751: code <= 4'b0000;
				752: code <= 4'bx101;
				753: code <= 4'b0001;
				754: code <= 4'b1000;
				755: code <= 4'bx111;
				756: code <= 4'b0000;
				757: code <= 4'bx111;
				758: code <= 4'b0010;
				759: code <= 4'b0001;
				760: code <= 4'b0001;
				761: code <= 4'bx011;
				762: code <= 4'bx100;
				763: code <= 4'b1001;
				764: code <= 4'b1001;
				765: code <= 4'b1001;
				766: code <= 4'b1001;
				767: code <= 4'b1001;
				768: code <= 4'b1001;
				769: code <= 4'b1000;
				770: code <= 4'bx011;
				771: code <= 4'bx111;
				772: code <= 4'b0010;
				773: code <= 4'b1001;
				774: code <= 4'bx111;
				775: code <= 4'b1000;
				776: code <= 4'b0000;
				777: code <= 4'bx100;
				778: code <= 4'b1001;
				779: code <= 4'b1001;
				780: code <= 4'bx101;
				781: code <= 4'b0001;
				782: code <= 4'b0000;
				783: code <= 4'bx101;
				784: code <= 4'b1001;
				785: code <= 4'bx111;
				786: code <= 4'bx011;
				787: code <= 4'b0001;
				788: code <= 4'bx111;
				789: code <= 4'bx011;
				790: code <= 4'b0010;
				791: code <= 4'b1000;
				792: code <= 4'b0001;
				793: code <= 4'bx110;
				794: code <= 4'b0000;
				795: code <= 4'b1001;
				796: code <= 4'bx110;
				797: code <= 4'bx011;
				798: code <= 4'b0001;
				799: code <= 4'b1000;
				800: code <= 4'bx101;
				801: code <= 4'b1001;
				802: code <= 4'bx101;
				803: code <= 4'b0000;
				804: code <= 4'b0010;
				805: code <= 4'bx100;
				806: code <= 4'bx100;
				807: code <= 4'bx101;
				808: code <= 4'b1001;
				809: code <= 4'bx100;
				810: code <= 4'bx101;
				811: code <= 4'bx101;
				812: code <= 4'bx011;
				813: code <= 4'bx100;
				814: code <= 4'bx110;
				815: code <= 4'b1001;
				816: code <= 4'b0000;
				817: code <= 4'b1000;
				818: code <= 4'bx011;
				819: code <= 4'b0000;
				820: code <= 4'b0010;
				821: code <= 4'bx110;
				822: code <= 4'bx100;
				823: code <= 4'b0010;
				824: code <= 4'bx101;
				825: code <= 4'b0010;
				826: code <= 4'b0010;
				827: code <= 4'bx011;
				828: code <= 4'b0000;
				829: code <= 4'b1000;
				830: code <= 4'b0010;
				831: code <= 4'bx101;
				832: code <= 4'bx011;
				833: code <= 4'bx011;
				834: code <= 4'bx100;
				835: code <= 4'bx100;
				836: code <= 4'bx110;
				837: code <= 4'b1000;
				838: code <= 4'bx101;
				839: code <= 4'b0000;
				840: code <= 4'bx011;
				841: code <= 4'bx101;
				842: code <= 4'b0010;
				843: code <= 4'bx110;
				844: code <= 4'b0001;
				845: code <= 4'b1001;
				846: code <= 4'bx011;
				847: code <= 4'b0001;
				848: code <= 4'b0001;
				849: code <= 4'b1000;
				850: code <= 4'b1000;
				851: code <= 4'b0001;
				852: code <= 4'bx111;
				853: code <= 4'b0001;
				854: code <= 4'b0000;
				855: code <= 4'b0001;
				856: code <= 4'b0000;
				857: code <= 4'b0000;
				858: code <= 4'b0000;
				859: code <= 4'bx011;
				860: code <= 4'b0001;
				861: code <= 4'bx011;
				862: code <= 4'bx111;
				863: code <= 4'b1000;
				864: code <= 4'bx011;
				865: code <= 4'b1000;
				866: code <= 4'bx111;
				867: code <= 4'bx101;
				868: code <= 4'b0010;
				869: code <= 4'b1000;
				870: code <= 4'b1000;
				871: code <= 4'bx110;
				872: code <= 4'bx101;
				873: code <= 4'b1000;
				874: code <= 4'bx111;
				875: code <= 4'bx101;
				876: code <= 4'bx011;
				877: code <= 4'bx011;
				878: code <= 4'b0010;
				879: code <= 4'b0000;
				880: code <= 4'b1000;
				881: code <= 4'bx011;
				882: code <= 4'b1000;
				883: code <= 4'b0001;
				884: code <= 4'bx100;
				885: code <= 4'b0010;
				886: code <= 4'b0000;
				887: code <= 4'bx110;
				888: code <= 4'b0001;
				889: code <= 4'bx111;
				890: code <= 4'b0001;
				891: code <= 4'bx111;
				892: code <= 4'bx111;
				893: code <= 4'bx110;
				894: code <= 4'bx110;
				895: code <= 4'b1001;
				896: code <= 4'b0001;
				897: code <= 4'bx100;
				898: code <= 4'bx111;
				899: code <= 4'bx011;
				900: code <= 4'b0000;
				901: code <= 4'bx011;
				902: code <= 4'bx101;
				903: code <= 4'b1001;
				904: code <= 4'b1000;
				905: code <= 4'b0010;
				906: code <= 4'bx101;
				907: code <= 4'bx011;
				908: code <= 4'bx100;
				909: code <= 4'b1001;
				910: code <= 4'b0000;
				911: code <= 4'bx100;
				912: code <= 4'b0010;
				913: code <= 4'b1000;
				914: code <= 4'bx111;
				915: code <= 4'bx101;
				916: code <= 4'bx101;
				917: code <= 4'bx100;
				918: code <= 4'bx110;
				919: code <= 4'b1000;
				920: code <= 4'bx111;
				921: code <= 4'bx011;
				922: code <= 4'b0001;
				923: code <= 4'b0001;
				924: code <= 4'bx101;
				925: code <= 4'b1001;
				926: code <= 4'bx101;
				927: code <= 4'bx110;
				928: code <= 4'b0010;
				929: code <= 4'b1000;
				930: code <= 4'bx110;
				931: code <= 4'bx011;
				932: code <= 4'b1000;
				933: code <= 4'b1000;
				934: code <= 4'b0010;
				935: code <= 4'bx011;
				936: code <= 4'bx101;
				937: code <= 4'bx011;
				938: code <= 4'bx111;
				939: code <= 4'b1000;
				940: code <= 4'bx111;
				941: code <= 4'bx101;
				942: code <= 4'b1001;
				943: code <= 4'bx011;
				944: code <= 4'bx111;
				945: code <= 4'bx101;
				946: code <= 4'b0001;
				947: code <= 4'b1001;
				948: code <= 4'bx101;
				949: code <= 4'bx111;
				950: code <= 4'bx111;
				951: code <= 4'b1000;
				952: code <= 4'b0001;
				953: code <= 4'b1000;
				954: code <= 4'bx101;
				955: code <= 4'bx111;
				956: code <= 4'bx111;
				957: code <= 4'b1000;
				958: code <= 4'b0000;
				959: code <= 4'bx101;
				960: code <= 4'bx011;
				961: code <= 4'b0010;
				962: code <= 4'b0001;
				963: code <= 4'bx111;
				964: code <= 4'b0001;
				965: code <= 4'b0010;
				966: code <= 4'b0010;
				967: code <= 4'bx110;
				968: code <= 4'b1000;
				969: code <= 4'b0000;
				970: code <= 4'bx110;
				971: code <= 4'bx110;
				972: code <= 4'b0001;
				973: code <= 4'bx011;
				974: code <= 4'b0000;
				975: code <= 4'b0000;
				976: code <= 4'b0001;
				977: code <= 4'b1001;
				978: code <= 4'b0010;
				979: code <= 4'bx111;
				980: code <= 4'b1000;
				981: code <= 4'bx111;
				982: code <= 4'bx110;
				983: code <= 4'bx110;
				984: code <= 4'b0001;
				985: code <= 4'b0001;
				986: code <= 4'b0001;
				987: code <= 4'b1001;
				988: code <= 4'bx101;
				989: code <= 4'b1001;
				990: code <= 4'b0000;
				991: code <= 4'b1001;
				992: code <= 4'b0010;
				993: code <= 4'b0001;
				994: code <= 4'bx110;
				995: code <= 4'bx100;
				996: code <= 4'b0010;
				997: code <= 4'b0000;
				998: code <= 4'b0001;
				999: code <= 4'b1001;
				1000: code <= 4'b1000;
				1001: code <= 4'b1001;
				1002: code <= 4'bx011;
				1003: code <= 4'b1000;
				1004: code <= 4'b0000;
				1005: code <= 4'b1001;
				1006: code <= 4'bx101;
				1007: code <= 4'b0010;
				1008: code <= 4'bx101;
				1009: code <= 4'bx111;
				1010: code <= 4'b0010;
				1011: code <= 4'b0000;
				1012: code <= 4'b0001;
				1013: code <= 4'b0000;
				1014: code <= 4'bx110;
				1015: code <= 4'bx101;
				1016: code <= 4'bx100;
				1017: code <= 4'b1000;
				1018: code <= 4'bx101;
				1019: code <= 4'b1000;
				1020: code <= 4'bx110;
				1021: code <= 4'bx011;
				1022: code <= 4'b0010;
				1023: code <= 4'bx111;
			endcase
			/* verilator lint_on CASEX */
		end
	end

	decoder decoder(.code(code), .segments(io_out));

endmodule

module jar_pi
(
	input  [7:0] io_in,
	output [7:0] io_out
);
	wire       clk      = io_in[0];
	wire       reset    = io_in[1];
//	wire       stream   = io_in[2];
//	wire [4:0] io_index = io_in[7:3];

	reg [9:0] index;
	//reg [7:0] led_out;
	reg [3:0] code;
	//assign io_out[7:0] = led_out;

	always @(posedge clk) begin
		if (reset) begin
//			index <= {io_index, index[9:5]};
			index <= 10'b0000000000;
		end
		else begin
//		else if (stream) begin
			index <= index + 1;
//		end

			case(index)
				10'd0: code <= 4'd3;
				10'd1: code <= 4'd10;
				10'd2: code <= 4'd1;
				10'd3: code <= 4'd4;
				10'd4: code <= 4'd1;
				10'd5: code <= 4'd5;
				10'd6: code <= 4'd9;
				10'd7: code <= 4'd2;
				10'd8: code <= 4'd6;
				10'd9: code <= 4'd5;
				10'd10: code <= 4'd3;
				10'd11: code <= 4'd5;
				10'd12: code <= 4'd8;
				10'd13: code <= 4'd9;
				10'd14: code <= 4'd7;
				10'd15: code <= 4'd9;
				10'd16: code <= 4'd3;
				10'd17: code <= 4'd2;
				10'd18: code <= 4'd3;
				10'd19: code <= 4'd8;
				10'd20: code <= 4'd4;
				10'd21: code <= 4'd6;
				10'd22: code <= 4'd2;
				10'd23: code <= 4'd6;
				10'd24: code <= 4'd4;
				10'd25: code <= 4'd3;
				10'd26: code <= 4'd3;
				10'd27: code <= 4'd8;
				10'd28: code <= 4'd3;
				10'd29: code <= 4'd2;
				10'd30: code <= 4'd7;
				10'd31: code <= 4'd9;
				10'd32: code <= 4'd5;
				10'd33: code <= 4'd0;
				10'd34: code <= 4'd2;
				10'd35: code <= 4'd8;
				10'd36: code <= 4'd8;
				10'd37: code <= 4'd4;
				10'd38: code <= 4'd1;
				10'd39: code <= 4'd9;
				10'd40: code <= 4'd7;
				10'd41: code <= 4'd1;
				10'd42: code <= 4'd6;
				10'd43: code <= 4'd9;
				10'd44: code <= 4'd3;
				10'd45: code <= 4'd9;
				10'd46: code <= 4'd9;
				10'd47: code <= 4'd3;
				10'd48: code <= 4'd7;
				10'd49: code <= 4'd5;
				10'd50: code <= 4'd1;
				10'd51: code <= 4'd0;
				10'd52: code <= 4'd5;
				10'd53: code <= 4'd8;
				10'd54: code <= 4'd2;
				10'd55: code <= 4'd0;
				10'd56: code <= 4'd9;
				10'd57: code <= 4'd7;
				10'd58: code <= 4'd4;
				10'd59: code <= 4'd9;
				10'd60: code <= 4'd4;
				10'd61: code <= 4'd4;
				10'd62: code <= 4'd5;
				10'd63: code <= 4'd9;
				10'd64: code <= 4'd2;
				10'd65: code <= 4'd3;
				10'd66: code <= 4'd0;
				10'd67: code <= 4'd7;
				10'd68: code <= 4'd8;
				10'd69: code <= 4'd1;
				10'd70: code <= 4'd6;
				10'd71: code <= 4'd4;
				10'd72: code <= 4'd0;
				10'd73: code <= 4'd6;
				10'd74: code <= 4'd2;
				10'd75: code <= 4'd8;
				10'd76: code <= 4'd6;
				10'd77: code <= 4'd2;
				10'd78: code <= 4'd0;
				10'd79: code <= 4'd8;
				10'd80: code <= 4'd9;
				10'd81: code <= 4'd9;
				10'd82: code <= 4'd8;
				10'd83: code <= 4'd6;
				10'd84: code <= 4'd2;
				10'd85: code <= 4'd8;
				10'd86: code <= 4'd0;
				10'd87: code <= 4'd3;
				10'd88: code <= 4'd4;
				10'd89: code <= 4'd8;
				10'd90: code <= 4'd2;
				10'd91: code <= 4'd5;
				10'd92: code <= 4'd3;
				10'd93: code <= 4'd4;
				10'd94: code <= 4'd2;
				10'd95: code <= 4'd1;
				10'd96: code <= 4'd1;
				10'd97: code <= 4'd7;
				10'd98: code <= 4'd0;
				10'd99: code <= 4'd6;
				10'd100: code <= 4'd7;
				10'd101: code <= 4'd9;
				10'd102: code <= 4'd8;
				10'd103: code <= 4'd2;
				10'd104: code <= 4'd1;
				10'd105: code <= 4'd4;
				10'd106: code <= 4'd8;
				10'd107: code <= 4'd0;
				10'd108: code <= 4'd8;
				10'd109: code <= 4'd6;
				10'd110: code <= 4'd5;
				10'd111: code <= 4'd1;
				10'd112: code <= 4'd3;
				10'd113: code <= 4'd2;
				10'd114: code <= 4'd8;
				10'd115: code <= 4'd2;
				10'd116: code <= 4'd3;
				10'd117: code <= 4'd0;
				10'd118: code <= 4'd6;
				10'd119: code <= 4'd6;
				10'd120: code <= 4'd4;
				10'd121: code <= 4'd7;
				10'd122: code <= 4'd0;
				10'd123: code <= 4'd9;
				10'd124: code <= 4'd3;
				10'd125: code <= 4'd8;
				10'd126: code <= 4'd4;
				10'd127: code <= 4'd4;
				10'd128: code <= 4'd6;
				10'd129: code <= 4'd0;
				10'd130: code <= 4'd9;
				10'd131: code <= 4'd5;
				10'd132: code <= 4'd5;
				10'd133: code <= 4'd0;
				10'd134: code <= 4'd5;
				10'd135: code <= 4'd8;
				10'd136: code <= 4'd2;
				10'd137: code <= 4'd2;
				10'd138: code <= 4'd3;
				10'd139: code <= 4'd1;
				10'd140: code <= 4'd7;
				10'd141: code <= 4'd2;
				10'd142: code <= 4'd5;
				10'd143: code <= 4'd3;
				10'd144: code <= 4'd5;
				10'd145: code <= 4'd9;
				10'd146: code <= 4'd4;
				10'd147: code <= 4'd0;
				10'd148: code <= 4'd8;
				10'd149: code <= 4'd1;
				10'd150: code <= 4'd2;
				10'd151: code <= 4'd8;
				10'd152: code <= 4'd4;
				10'd153: code <= 4'd8;
				10'd154: code <= 4'd1;
				10'd155: code <= 4'd1;
				10'd156: code <= 4'd1;
				10'd157: code <= 4'd7;
				10'd158: code <= 4'd4;
				10'd159: code <= 4'd5;
				10'd160: code <= 4'd0;
				10'd161: code <= 4'd2;
				10'd162: code <= 4'd8;
				10'd163: code <= 4'd4;
				10'd164: code <= 4'd1;
				10'd165: code <= 4'd0;
				10'd166: code <= 4'd2;
				10'd167: code <= 4'd7;
				10'd168: code <= 4'd0;
				10'd169: code <= 4'd1;
				10'd170: code <= 4'd9;
				10'd171: code <= 4'd3;
				10'd172: code <= 4'd8;
				10'd173: code <= 4'd5;
				10'd174: code <= 4'd2;
				10'd175: code <= 4'd1;
				10'd176: code <= 4'd1;
				10'd177: code <= 4'd0;
				10'd178: code <= 4'd5;
				10'd179: code <= 4'd5;
				10'd180: code <= 4'd5;
				10'd181: code <= 4'd9;
				10'd182: code <= 4'd6;
				10'd183: code <= 4'd4;
				10'd184: code <= 4'd4;
				10'd185: code <= 4'd6;
				10'd186: code <= 4'd2;
				10'd187: code <= 4'd2;
				10'd188: code <= 4'd9;
				10'd189: code <= 4'd4;
				10'd190: code <= 4'd8;
				10'd191: code <= 4'd9;
				10'd192: code <= 4'd5;
				10'd193: code <= 4'd4;
				10'd194: code <= 4'd9;
				10'd195: code <= 4'd3;
				10'd196: code <= 4'd0;
				10'd197: code <= 4'd3;
				10'd198: code <= 4'd8;
				10'd199: code <= 4'd1;
				10'd200: code <= 4'd9;
				10'd201: code <= 4'd6;
				10'd202: code <= 4'd4;
				10'd203: code <= 4'd4;
				10'd204: code <= 4'd2;
				10'd205: code <= 4'd8;
				10'd206: code <= 4'd8;
				10'd207: code <= 4'd1;
				10'd208: code <= 4'd0;
				10'd209: code <= 4'd9;
				10'd210: code <= 4'd7;
				10'd211: code <= 4'd5;
				10'd212: code <= 4'd6;
				10'd213: code <= 4'd6;
				10'd214: code <= 4'd5;
				10'd215: code <= 4'd9;
				10'd216: code <= 4'd3;
				10'd217: code <= 4'd3;
				10'd218: code <= 4'd4;
				10'd219: code <= 4'd4;
				10'd220: code <= 4'd6;
				10'd221: code <= 4'd1;
				10'd222: code <= 4'd2;
				10'd223: code <= 4'd8;
				10'd224: code <= 4'd4;
				10'd225: code <= 4'd7;
				10'd226: code <= 4'd5;
				10'd227: code <= 4'd6;
				10'd228: code <= 4'd4;
				10'd229: code <= 4'd8;
				10'd230: code <= 4'd2;
				10'd231: code <= 4'd3;
				10'd232: code <= 4'd3;
				10'd233: code <= 4'd7;
				10'd234: code <= 4'd8;
				10'd235: code <= 4'd6;
				10'd236: code <= 4'd7;
				10'd237: code <= 4'd8;
				10'd238: code <= 4'd3;
				10'd239: code <= 4'd1;
				10'd240: code <= 4'd6;
				10'd241: code <= 4'd5;
				10'd242: code <= 4'd2;
				10'd243: code <= 4'd7;
				10'd244: code <= 4'd1;
				10'd245: code <= 4'd2;
				10'd246: code <= 4'd0;
				10'd247: code <= 4'd1;
				10'd248: code <= 4'd9;
				10'd249: code <= 4'd0;
				10'd250: code <= 4'd9;
				10'd251: code <= 4'd1;
				10'd252: code <= 4'd4;
				10'd253: code <= 4'd5;
				10'd254: code <= 4'd6;
				10'd255: code <= 4'd4;
				10'd256: code <= 4'd8;
				10'd257: code <= 4'd5;
				10'd258: code <= 4'd6;
				10'd259: code <= 4'd6;
				10'd260: code <= 4'd9;
				10'd261: code <= 4'd2;
				10'd262: code <= 4'd3;
				10'd263: code <= 4'd4;
				10'd264: code <= 4'd6;
				10'd265: code <= 4'd0;
				10'd266: code <= 4'd3;
				10'd267: code <= 4'd4;
				10'd268: code <= 4'd8;
				10'd269: code <= 4'd6;
				10'd270: code <= 4'd1;
				10'd271: code <= 4'd0;
				10'd272: code <= 4'd4;
				10'd273: code <= 4'd5;
				10'd274: code <= 4'd4;
				10'd275: code <= 4'd3;
				10'd276: code <= 4'd2;
				10'd277: code <= 4'd6;
				10'd278: code <= 4'd6;
				10'd279: code <= 4'd4;
				10'd280: code <= 4'd8;
				10'd281: code <= 4'd2;
				10'd282: code <= 4'd1;
				10'd283: code <= 4'd3;
				10'd284: code <= 4'd3;
				10'd285: code <= 4'd9;
				10'd286: code <= 4'd3;
				10'd287: code <= 4'd6;
				10'd288: code <= 4'd0;
				10'd289: code <= 4'd7;
				10'd290: code <= 4'd2;
				10'd291: code <= 4'd6;
				10'd292: code <= 4'd0;
				10'd293: code <= 4'd2;
				10'd294: code <= 4'd4;
				10'd295: code <= 4'd9;
				10'd296: code <= 4'd1;
				10'd297: code <= 4'd4;
				10'd298: code <= 4'd1;
				10'd299: code <= 4'd2;
				10'd300: code <= 4'd7;
				10'd301: code <= 4'd3;
				10'd302: code <= 4'd7;
				10'd303: code <= 4'd2;
				10'd304: code <= 4'd4;
				10'd305: code <= 4'd5;
				10'd306: code <= 4'd8;
				10'd307: code <= 4'd7;
				10'd308: code <= 4'd0;
				10'd309: code <= 4'd0;
				10'd310: code <= 4'd6;
				10'd311: code <= 4'd6;
				10'd312: code <= 4'd0;
				10'd313: code <= 4'd6;
				10'd314: code <= 4'd3;
				10'd315: code <= 4'd1;
				10'd316: code <= 4'd5;
				10'd317: code <= 4'd5;
				10'd318: code <= 4'd8;
				10'd319: code <= 4'd8;
				10'd320: code <= 4'd1;
				10'd321: code <= 4'd7;
				10'd322: code <= 4'd4;
				10'd323: code <= 4'd8;
				10'd324: code <= 4'd8;
				10'd325: code <= 4'd1;
				10'd326: code <= 4'd5;
				10'd327: code <= 4'd2;
				10'd328: code <= 4'd0;
				10'd329: code <= 4'd9;
				10'd330: code <= 4'd2;
				10'd331: code <= 4'd0;
				10'd332: code <= 4'd9;
				10'd333: code <= 4'd6;
				10'd334: code <= 4'd2;
				10'd335: code <= 4'd8;
				10'd336: code <= 4'd2;
				10'd337: code <= 4'd9;
				10'd338: code <= 4'd2;
				10'd339: code <= 4'd5;
				10'd340: code <= 4'd4;
				10'd341: code <= 4'd0;
				10'd342: code <= 4'd9;
				10'd343: code <= 4'd1;
				10'd344: code <= 4'd7;
				10'd345: code <= 4'd1;
				10'd346: code <= 4'd5;
				10'd347: code <= 4'd3;
				10'd348: code <= 4'd6;
				10'd349: code <= 4'd4;
				10'd350: code <= 4'd3;
				10'd351: code <= 4'd6;
				10'd352: code <= 4'd7;
				10'd353: code <= 4'd8;
				10'd354: code <= 4'd9;
				10'd355: code <= 4'd2;
				10'd356: code <= 4'd5;
				10'd357: code <= 4'd9;
				10'd358: code <= 4'd0;
				10'd359: code <= 4'd3;
				10'd360: code <= 4'd6;
				10'd361: code <= 4'd0;
				10'd362: code <= 4'd0;
				10'd363: code <= 4'd1;
				10'd364: code <= 4'd1;
				10'd365: code <= 4'd3;
				10'd366: code <= 4'd3;
				10'd367: code <= 4'd0;
				10'd368: code <= 4'd5;
				10'd369: code <= 4'd3;
				10'd370: code <= 4'd0;
				10'd371: code <= 4'd5;
				10'd372: code <= 4'd4;
				10'd373: code <= 4'd8;
				10'd374: code <= 4'd8;
				10'd375: code <= 4'd2;
				10'd376: code <= 4'd0;
				10'd377: code <= 4'd4;
				10'd378: code <= 4'd6;
				10'd379: code <= 4'd6;
				10'd380: code <= 4'd5;
				10'd381: code <= 4'd2;
				10'd382: code <= 4'd1;
				10'd383: code <= 4'd3;
				10'd384: code <= 4'd8;
				10'd385: code <= 4'd4;
				10'd386: code <= 4'd1;
				10'd387: code <= 4'd4;
				10'd388: code <= 4'd6;
				10'd389: code <= 4'd9;
				10'd390: code <= 4'd5;
				10'd391: code <= 4'd1;
				10'd392: code <= 4'd9;
				10'd393: code <= 4'd4;
				10'd394: code <= 4'd1;
				10'd395: code <= 4'd5;
				10'd396: code <= 4'd1;
				10'd397: code <= 4'd1;
				10'd398: code <= 4'd6;
				10'd399: code <= 4'd0;
				10'd400: code <= 4'd9;
				10'd401: code <= 4'd4;
				10'd402: code <= 4'd3;
				10'd403: code <= 4'd3;
				10'd404: code <= 4'd0;
				10'd405: code <= 4'd5;
				10'd406: code <= 4'd7;
				10'd407: code <= 4'd2;
				10'd408: code <= 4'd7;
				10'd409: code <= 4'd0;
				10'd410: code <= 4'd3;
				10'd411: code <= 4'd6;
				10'd412: code <= 4'd5;
				10'd413: code <= 4'd7;
				10'd414: code <= 4'd5;
				10'd415: code <= 4'd9;
				10'd416: code <= 4'd5;
				10'd417: code <= 4'd9;
				10'd418: code <= 4'd1;
				10'd419: code <= 4'd9;
				10'd420: code <= 4'd5;
				10'd421: code <= 4'd3;
				10'd422: code <= 4'd0;
				10'd423: code <= 4'd9;
				10'd424: code <= 4'd2;
				10'd425: code <= 4'd1;
				10'd426: code <= 4'd8;
				10'd427: code <= 4'd6;
				10'd428: code <= 4'd1;
				10'd429: code <= 4'd1;
				10'd430: code <= 4'd7;
				10'd431: code <= 4'd3;
				10'd432: code <= 4'd8;
				10'd433: code <= 4'd1;
				10'd434: code <= 4'd9;
				10'd435: code <= 4'd3;
				10'd436: code <= 4'd2;
				10'd437: code <= 4'd6;
				10'd438: code <= 4'd1;
				10'd439: code <= 4'd1;
				10'd440: code <= 4'd7;
				10'd441: code <= 4'd9;
				10'd442: code <= 4'd3;
				10'd443: code <= 4'd1;
				10'd444: code <= 4'd0;
				10'd445: code <= 4'd5;
				10'd446: code <= 4'd1;
				10'd447: code <= 4'd1;
				10'd448: code <= 4'd8;
				10'd449: code <= 4'd5;
				10'd450: code <= 4'd4;
				10'd451: code <= 4'd8;
				10'd452: code <= 4'd0;
				10'd453: code <= 4'd7;
				10'd454: code <= 4'd4;
				10'd455: code <= 4'd4;
				10'd456: code <= 4'd6;
				10'd457: code <= 4'd2;
				10'd458: code <= 4'd3;
				10'd459: code <= 4'd7;
				10'd460: code <= 4'd9;
				10'd461: code <= 4'd9;
				10'd462: code <= 4'd6;
				10'd463: code <= 4'd2;
				10'd464: code <= 4'd7;
				10'd465: code <= 4'd4;
				10'd466: code <= 4'd9;
				10'd467: code <= 4'd5;
				10'd468: code <= 4'd6;
				10'd469: code <= 4'd7;
				10'd470: code <= 4'd3;
				10'd471: code <= 4'd5;
				10'd472: code <= 4'd1;
				10'd473: code <= 4'd8;
				10'd474: code <= 4'd8;
				10'd475: code <= 4'd5;
				10'd476: code <= 4'd7;
				10'd477: code <= 4'd5;
				10'd478: code <= 4'd2;
				10'd479: code <= 4'd7;
				10'd480: code <= 4'd2;
				10'd481: code <= 4'd4;
				10'd482: code <= 4'd8;
				10'd483: code <= 4'd9;
				10'd484: code <= 4'd1;
				10'd485: code <= 4'd2;
				10'd486: code <= 4'd2;
				10'd487: code <= 4'd7;
				10'd488: code <= 4'd9;
				10'd489: code <= 4'd3;
				10'd490: code <= 4'd8;
				10'd491: code <= 4'd1;
				10'd492: code <= 4'd8;
				10'd493: code <= 4'd3;
				10'd494: code <= 4'd0;
				10'd495: code <= 4'd1;
				10'd496: code <= 4'd1;
				10'd497: code <= 4'd9;
				10'd498: code <= 4'd4;
				10'd499: code <= 4'd9;
				10'd500: code <= 4'd1;
				10'd501: code <= 4'd2;
				10'd502: code <= 4'd9;
				10'd503: code <= 4'd8;
				10'd504: code <= 4'd3;
				10'd505: code <= 4'd3;
				10'd506: code <= 4'd6;
				10'd507: code <= 4'd7;
				10'd508: code <= 4'd3;
				10'd509: code <= 4'd3;
				10'd510: code <= 4'd6;
				10'd511: code <= 4'd2;
				10'd512: code <= 4'd4;
				10'd513: code <= 4'd4;
				10'd514: code <= 4'd0;
				10'd515: code <= 4'd6;
				10'd516: code <= 4'd5;
				10'd517: code <= 4'd6;
				10'd518: code <= 4'd6;
				10'd519: code <= 4'd4;
				10'd520: code <= 4'd3;
				10'd521: code <= 4'd0;
				10'd522: code <= 4'd8;
				10'd523: code <= 4'd6;
				10'd524: code <= 4'd0;
				10'd525: code <= 4'd2;
				10'd526: code <= 4'd1;
				10'd527: code <= 4'd3;
				10'd528: code <= 4'd9;
				10'd529: code <= 4'd4;
				10'd530: code <= 4'd9;
				10'd531: code <= 4'd4;
				10'd532: code <= 4'd6;
				10'd533: code <= 4'd3;
				10'd534: code <= 4'd9;
				10'd535: code <= 4'd5;
				10'd536: code <= 4'd2;
				10'd537: code <= 4'd2;
				10'd538: code <= 4'd4;
				10'd539: code <= 4'd7;
				10'd540: code <= 4'd3;
				10'd541: code <= 4'd7;
				10'd542: code <= 4'd1;
				10'd543: code <= 4'd9;
				10'd544: code <= 4'd0;
				10'd545: code <= 4'd7;
				10'd546: code <= 4'd0;
				10'd547: code <= 4'd2;
				10'd548: code <= 4'd1;
				10'd549: code <= 4'd7;
				10'd550: code <= 4'd9;
				10'd551: code <= 4'd8;
				10'd552: code <= 4'd6;
				10'd553: code <= 4'd0;
				10'd554: code <= 4'd9;
				10'd555: code <= 4'd4;
				10'd556: code <= 4'd3;
				10'd557: code <= 4'd7;
				10'd558: code <= 4'd0;
				10'd559: code <= 4'd2;
				10'd560: code <= 4'd7;
				10'd561: code <= 4'd7;
				10'd562: code <= 4'd0;
				10'd563: code <= 4'd5;
				10'd564: code <= 4'd3;
				10'd565: code <= 4'd9;
				10'd566: code <= 4'd2;
				10'd567: code <= 4'd1;
				10'd568: code <= 4'd7;
				10'd569: code <= 4'd1;
				10'd570: code <= 4'd7;
				10'd571: code <= 4'd6;
				10'd572: code <= 4'd2;
				10'd573: code <= 4'd9;
				10'd574: code <= 4'd3;
				10'd575: code <= 4'd1;
				10'd576: code <= 4'd7;
				10'd577: code <= 4'd6;
				10'd578: code <= 4'd7;
				10'd579: code <= 4'd5;
				10'd580: code <= 4'd2;
				10'd581: code <= 4'd3;
				10'd582: code <= 4'd8;
				10'd583: code <= 4'd4;
				10'd584: code <= 4'd6;
				10'd585: code <= 4'd7;
				10'd586: code <= 4'd4;
				10'd587: code <= 4'd8;
				10'd588: code <= 4'd1;
				10'd589: code <= 4'd8;
				10'd590: code <= 4'd4;
				10'd591: code <= 4'd6;
				10'd592: code <= 4'd7;
				10'd593: code <= 4'd6;
				10'd594: code <= 4'd6;
				10'd595: code <= 4'd9;
				10'd596: code <= 4'd4;
				10'd597: code <= 4'd0;
				10'd598: code <= 4'd5;
				10'd599: code <= 4'd1;
				10'd600: code <= 4'd3;
				10'd601: code <= 4'd2;
				10'd602: code <= 4'd0;
				10'd603: code <= 4'd0;
				10'd604: code <= 4'd0;
				10'd605: code <= 4'd5;
				10'd606: code <= 4'd6;
				10'd607: code <= 4'd8;
				10'd608: code <= 4'd1;
				10'd609: code <= 4'd2;
				10'd610: code <= 4'd7;
				10'd611: code <= 4'd1;
				10'd612: code <= 4'd4;
				10'd613: code <= 4'd5;
				10'd614: code <= 4'd2;
				10'd615: code <= 4'd6;
				10'd616: code <= 4'd3;
				10'd617: code <= 4'd5;
				10'd618: code <= 4'd6;
				10'd619: code <= 4'd0;
				10'd620: code <= 4'd8;
				10'd621: code <= 4'd2;
				10'd622: code <= 4'd7;
				10'd623: code <= 4'd7;
				10'd624: code <= 4'd8;
				10'd625: code <= 4'd5;
				10'd626: code <= 4'd7;
				10'd627: code <= 4'd7;
				10'd628: code <= 4'd1;
				10'd629: code <= 4'd3;
				10'd630: code <= 4'd4;
				10'd631: code <= 4'd2;
				10'd632: code <= 4'd7;
				10'd633: code <= 4'd5;
				10'd634: code <= 4'd7;
				10'd635: code <= 4'd7;
				10'd636: code <= 4'd8;
				10'd637: code <= 4'd9;
				10'd638: code <= 4'd6;
				10'd639: code <= 4'd0;
				10'd640: code <= 4'd9;
				10'd641: code <= 4'd1;
				10'd642: code <= 4'd7;
				10'd643: code <= 4'd3;
				10'd644: code <= 4'd6;
				10'd645: code <= 4'd3;
				10'd646: code <= 4'd7;
				10'd647: code <= 4'd1;
				10'd648: code <= 4'd7;
				10'd649: code <= 4'd8;
				10'd650: code <= 4'd7;
				10'd651: code <= 4'd2;
				10'd652: code <= 4'd1;
				10'd653: code <= 4'd4;
				10'd654: code <= 4'd6;
				10'd655: code <= 4'd8;
				10'd656: code <= 4'd4;
				10'd657: code <= 4'd4;
				10'd658: code <= 4'd0;
				10'd659: code <= 4'd9;
				10'd660: code <= 4'd0;
				10'd661: code <= 4'd1;
				10'd662: code <= 4'd2;
				10'd663: code <= 4'd2;
				10'd664: code <= 4'd4;
				10'd665: code <= 4'd9;
				10'd666: code <= 4'd5;
				10'd667: code <= 4'd3;
				10'd668: code <= 4'd4;
				10'd669: code <= 4'd3;
				10'd670: code <= 4'd0;
				10'd671: code <= 4'd1;
				10'd672: code <= 4'd4;
				10'd673: code <= 4'd6;
				10'd674: code <= 4'd5;
				10'd675: code <= 4'd4;
				10'd676: code <= 4'd9;
				10'd677: code <= 4'd5;
				10'd678: code <= 4'd8;
				10'd679: code <= 4'd5;
				10'd680: code <= 4'd3;
				10'd681: code <= 4'd7;
				10'd682: code <= 4'd1;
				10'd683: code <= 4'd0;
				10'd684: code <= 4'd5;
				10'd685: code <= 4'd0;
				10'd686: code <= 4'd7;
				10'd687: code <= 4'd9;
				10'd688: code <= 4'd2;
				10'd689: code <= 4'd2;
				10'd690: code <= 4'd7;
				10'd691: code <= 4'd9;
				10'd692: code <= 4'd6;
				10'd693: code <= 4'd8;
				10'd694: code <= 4'd9;
				10'd695: code <= 4'd2;
				10'd696: code <= 4'd5;
				10'd697: code <= 4'd8;
				10'd698: code <= 4'd9;
				10'd699: code <= 4'd2;
				10'd700: code <= 4'd3;
				10'd701: code <= 4'd5;
				10'd702: code <= 4'd4;
				10'd703: code <= 4'd2;
				10'd704: code <= 4'd0;
				10'd705: code <= 4'd1;
				10'd706: code <= 4'd9;
				10'd707: code <= 4'd9;
				10'd708: code <= 4'd5;
				10'd709: code <= 4'd6;
				10'd710: code <= 4'd1;
				10'd711: code <= 4'd1;
				10'd712: code <= 4'd2;
				10'd713: code <= 4'd1;
				10'd714: code <= 4'd2;
				10'd715: code <= 4'd9;
				10'd716: code <= 4'd0;
				10'd717: code <= 4'd2;
				10'd718: code <= 4'd1;
				10'd719: code <= 4'd9;
				10'd720: code <= 4'd6;
				10'd721: code <= 4'd0;
				10'd722: code <= 4'd8;
				10'd723: code <= 4'd6;
				10'd724: code <= 4'd4;
				10'd725: code <= 4'd0;
				10'd726: code <= 4'd3;
				10'd727: code <= 4'd4;
				10'd728: code <= 4'd4;
				10'd729: code <= 4'd1;
				10'd730: code <= 4'd8;
				10'd731: code <= 4'd1;
				10'd732: code <= 4'd5;
				10'd733: code <= 4'd9;
				10'd734: code <= 4'd8;
				10'd735: code <= 4'd1;
				10'd736: code <= 4'd3;
				10'd737: code <= 4'd6;
				10'd738: code <= 4'd2;
				10'd739: code <= 4'd9;
				10'd740: code <= 4'd7;
				10'd741: code <= 4'd7;
				10'd742: code <= 4'd4;
				10'd743: code <= 4'd7;
				10'd744: code <= 4'd7;
				10'd745: code <= 4'd1;
				10'd746: code <= 4'd3;
				10'd747: code <= 4'd0;
				10'd748: code <= 4'd9;
				10'd749: code <= 4'd9;
				10'd750: code <= 4'd6;
				10'd751: code <= 4'd0;
				10'd752: code <= 4'd5;
				10'd753: code <= 4'd1;
				10'd754: code <= 4'd8;
				10'd755: code <= 4'd7;
				10'd756: code <= 4'd0;
				10'd757: code <= 4'd7;
				10'd758: code <= 4'd2;
				10'd759: code <= 4'd1;
				10'd760: code <= 4'd1;
				10'd761: code <= 4'd3;
				10'd762: code <= 4'd4;
				10'd763: code <= 4'd9;
				10'd764: code <= 4'd9;
				10'd765: code <= 4'd9;
				10'd766: code <= 4'd9;
				10'd767: code <= 4'd9;
				10'd768: code <= 4'd9;
				10'd769: code <= 4'd8;
				10'd770: code <= 4'd3;
				10'd771: code <= 4'd7;
				10'd772: code <= 4'd2;
				10'd773: code <= 4'd9;
				10'd774: code <= 4'd7;
				10'd775: code <= 4'd8;
				10'd776: code <= 4'd0;
				10'd777: code <= 4'd4;
				10'd778: code <= 4'd9;
				10'd779: code <= 4'd9;
				10'd780: code <= 4'd5;
				10'd781: code <= 4'd1;
				10'd782: code <= 4'd0;
				10'd783: code <= 4'd5;
				10'd784: code <= 4'd9;
				10'd785: code <= 4'd7;
				10'd786: code <= 4'd3;
				10'd787: code <= 4'd1;
				10'd788: code <= 4'd7;
				10'd789: code <= 4'd3;
				10'd790: code <= 4'd2;
				10'd791: code <= 4'd8;
				10'd792: code <= 4'd1;
				10'd793: code <= 4'd6;
				10'd794: code <= 4'd0;
				10'd795: code <= 4'd9;
				10'd796: code <= 4'd6;
				10'd797: code <= 4'd3;
				10'd798: code <= 4'd1;
				10'd799: code <= 4'd8;
				10'd800: code <= 4'd5;
				10'd801: code <= 4'd9;
				10'd802: code <= 4'd5;
				10'd803: code <= 4'd0;
				10'd804: code <= 4'd2;
				10'd805: code <= 4'd4;
				10'd806: code <= 4'd4;
				10'd807: code <= 4'd5;
				10'd808: code <= 4'd9;
				10'd809: code <= 4'd4;
				10'd810: code <= 4'd5;
				10'd811: code <= 4'd5;
				10'd812: code <= 4'd3;
				10'd813: code <= 4'd4;
				10'd814: code <= 4'd6;
				10'd815: code <= 4'd9;
				10'd816: code <= 4'd0;
				10'd817: code <= 4'd8;
				10'd818: code <= 4'd3;
				10'd819: code <= 4'd0;
				10'd820: code <= 4'd2;
				10'd821: code <= 4'd6;
				10'd822: code <= 4'd4;
				10'd823: code <= 4'd2;
				10'd824: code <= 4'd5;
				10'd825: code <= 4'd2;
				10'd826: code <= 4'd2;
				10'd827: code <= 4'd3;
				10'd828: code <= 4'd0;
				10'd829: code <= 4'd8;
				10'd830: code <= 4'd2;
				10'd831: code <= 4'd5;
				10'd832: code <= 4'd3;
				10'd833: code <= 4'd3;
				10'd834: code <= 4'd4;
				10'd835: code <= 4'd4;
				10'd836: code <= 4'd6;
				10'd837: code <= 4'd8;
				10'd838: code <= 4'd5;
				10'd839: code <= 4'd0;
				10'd840: code <= 4'd3;
				10'd841: code <= 4'd5;
				10'd842: code <= 4'd2;
				10'd843: code <= 4'd6;
				10'd844: code <= 4'd1;
				10'd845: code <= 4'd9;
				10'd846: code <= 4'd3;
				10'd847: code <= 4'd1;
				10'd848: code <= 4'd1;
				10'd849: code <= 4'd8;
				10'd850: code <= 4'd8;
				10'd851: code <= 4'd1;
				10'd852: code <= 4'd7;
				10'd853: code <= 4'd1;
				10'd854: code <= 4'd0;
				10'd855: code <= 4'd1;
				10'd856: code <= 4'd0;
				10'd857: code <= 4'd0;
				10'd858: code <= 4'd0;
				10'd859: code <= 4'd3;
				10'd860: code <= 4'd1;
				10'd861: code <= 4'd3;
				10'd862: code <= 4'd7;
				10'd863: code <= 4'd8;
				10'd864: code <= 4'd3;
				10'd865: code <= 4'd8;
				10'd866: code <= 4'd7;
				10'd867: code <= 4'd5;
				10'd868: code <= 4'd2;
				10'd869: code <= 4'd8;
				10'd870: code <= 4'd8;
				10'd871: code <= 4'd6;
				10'd872: code <= 4'd5;
				10'd873: code <= 4'd8;
				10'd874: code <= 4'd7;
				10'd875: code <= 4'd5;
				10'd876: code <= 4'd3;
				10'd877: code <= 4'd3;
				10'd878: code <= 4'd2;
				10'd879: code <= 4'd0;
				10'd880: code <= 4'd8;
				10'd881: code <= 4'd3;
				10'd882: code <= 4'd8;
				10'd883: code <= 4'd1;
				10'd884: code <= 4'd4;
				10'd885: code <= 4'd2;
				10'd886: code <= 4'd0;
				10'd887: code <= 4'd6;
				10'd888: code <= 4'd1;
				10'd889: code <= 4'd7;
				10'd890: code <= 4'd1;
				10'd891: code <= 4'd7;
				10'd892: code <= 4'd7;
				10'd893: code <= 4'd6;
				10'd894: code <= 4'd6;
				10'd895: code <= 4'd9;
				10'd896: code <= 4'd1;
				10'd897: code <= 4'd4;
				10'd898: code <= 4'd7;
				10'd899: code <= 4'd3;
				10'd900: code <= 4'd0;
				10'd901: code <= 4'd3;
				10'd902: code <= 4'd5;
				10'd903: code <= 4'd9;
				10'd904: code <= 4'd8;
				10'd905: code <= 4'd2;
				10'd906: code <= 4'd5;
				10'd907: code <= 4'd3;
				10'd908: code <= 4'd4;
				10'd909: code <= 4'd9;
				10'd910: code <= 4'd0;
				10'd911: code <= 4'd4;
				10'd912: code <= 4'd2;
				10'd913: code <= 4'd8;
				10'd914: code <= 4'd7;
				10'd915: code <= 4'd5;
				10'd916: code <= 4'd5;
				10'd917: code <= 4'd4;
				10'd918: code <= 4'd6;
				10'd919: code <= 4'd8;
				10'd920: code <= 4'd7;
				10'd921: code <= 4'd3;
				10'd922: code <= 4'd1;
				10'd923: code <= 4'd1;
				10'd924: code <= 4'd5;
				10'd925: code <= 4'd9;
				10'd926: code <= 4'd5;
				10'd927: code <= 4'd6;
				10'd928: code <= 4'd2;
				10'd929: code <= 4'd8;
				10'd930: code <= 4'd6;
				10'd931: code <= 4'd3;
				10'd932: code <= 4'd8;
				10'd933: code <= 4'd8;
				10'd934: code <= 4'd2;
				10'd935: code <= 4'd3;
				10'd936: code <= 4'd5;
				10'd937: code <= 4'd3;
				10'd938: code <= 4'd7;
				10'd939: code <= 4'd8;
				10'd940: code <= 4'd7;
				10'd941: code <= 4'd5;
				10'd942: code <= 4'd9;
				10'd943: code <= 4'd3;
				10'd944: code <= 4'd7;
				10'd945: code <= 4'd5;
				10'd946: code <= 4'd1;
				10'd947: code <= 4'd9;
				10'd948: code <= 4'd5;
				10'd949: code <= 4'd7;
				10'd950: code <= 4'd7;
				10'd951: code <= 4'd8;
				10'd952: code <= 4'd1;
				10'd953: code <= 4'd8;
				10'd954: code <= 4'd5;
				10'd955: code <= 4'd7;
				10'd956: code <= 4'd7;
				10'd957: code <= 4'd8;
				10'd958: code <= 4'd0;
				10'd959: code <= 4'd5;
				10'd960: code <= 4'd3;
				10'd961: code <= 4'd2;
				10'd962: code <= 4'd1;
				10'd963: code <= 4'd7;
				10'd964: code <= 4'd1;
				10'd965: code <= 4'd2;
				10'd966: code <= 4'd2;
				10'd967: code <= 4'd6;
				10'd968: code <= 4'd8;
				10'd969: code <= 4'd0;
				10'd970: code <= 4'd6;
				10'd971: code <= 4'd6;
				10'd972: code <= 4'd1;
				10'd973: code <= 4'd3;
				10'd974: code <= 4'd0;
				10'd975: code <= 4'd0;
				10'd976: code <= 4'd1;
				10'd977: code <= 4'd9;
				10'd978: code <= 4'd2;
				10'd979: code <= 4'd7;
				10'd980: code <= 4'd8;
				10'd981: code <= 4'd7;
				10'd982: code <= 4'd6;
				10'd983: code <= 4'd6;
				10'd984: code <= 4'd1;
				10'd985: code <= 4'd1;
				10'd986: code <= 4'd1;
				10'd987: code <= 4'd9;
				10'd988: code <= 4'd5;
				10'd989: code <= 4'd9;
				10'd990: code <= 4'd0;
				10'd991: code <= 4'd9;
				10'd992: code <= 4'd2;
				10'd993: code <= 4'd1;
				10'd994: code <= 4'd6;
				10'd995: code <= 4'd4;
				10'd996: code <= 4'd2;
				10'd997: code <= 4'd0;
				10'd998: code <= 4'd1;
				10'd999: code <= 4'd9;
				10'd1000: code <= 4'd8;
				10'd1001: code <= 4'd9;
				10'd1002: code <= 4'd3;
				10'd1003: code <= 4'd8;
				10'd1004: code <= 4'd0;
				10'd1005: code <= 4'd9;
				10'd1006: code <= 4'd5;
				10'd1007: code <= 4'd2;
				10'd1008: code <= 4'd5;
				10'd1009: code <= 4'd7;
				10'd1010: code <= 4'd2;
				10'd1011: code <= 4'd0;
				10'd1012: code <= 4'd1;
				10'd1013: code <= 4'd0;
				10'd1014: code <= 4'd6;
				10'd1015: code <= 4'd5;
				10'd1016: code <= 4'd4;
				10'd1017: code <= 4'd8;
				10'd1018: code <= 4'd5;
				10'd1019: code <= 4'd8;
				10'd1020: code <= 4'd6;
				10'd1021: code <= 4'd3;
				10'd1022: code <= 4'd2;
				10'd1023: code <= 4'd7;
			endcase
		end
	end

	decoder decoder(.code(code), .segments(io_out));

endmodule

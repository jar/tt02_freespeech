module jar_pi
(
	input  [7:0] io_in,
	output [7:0] io_out
);
	wire       clk      = io_in[0];
	wire       reset    = io_in[1];
//	wire       stream   = io_in[2];
//	wire [4:0] io_index = io_in[7:3];

	reg [9:0] index;
	//reg [7:0] led_out;
	wire [3:0] code;
	//assign io_out[7:0] = led_out;

	wire j = index[9];
	wire i = index[8];
	wire h = index[7];
	wire g = index[6];
	wire f = index[5];
	wire e = index[4];
	wire d = index[3];
	wire c = index[2];
	wire b = index[1];
	wire a = index[0];

	always @(posedge clk) begin
		if (reset) begin
//			index <= {io_index, index[9:5]};
			index <= 10'b0000000000;
		end
		else begin
//		else if (stream) begin
			index <= index + 1;
//		end

code[3]<=j?((!i&!h&!g&f&!e&!d&c&b&!a)|(i&h&g&!f&e&d&b&a)|(!h&!g&!f&e&d&!c&b&a)|(!i&!h&!g&!f&e&!d&b&!a)|(!i&h&!g&e&d&!c&b&!a)|(!h&!g&f&!e&!d&!c&!b&a)|(!i&g&!f&!e&d&b&a)|(!i&!h&g&!f&d&c&a)|(!i&!h&!f&!d&c&b&!a)|(!h&g&f&e&!d&!c&!a)|(h&!g&!f&!e&d&c&a)|(i&!h&f&!e&!d&c&b)|(h&g&f&d&c&!b&a)|(h&!g&e&!d&!c&b&a)|(i&h&!g&!e&!d&b&a)|(!i&h&g&f&e&d&c)|(i&!h&!g&!e&d&b&a)|(!i&h&!g&!f&!e&!c&!a)|(!i&h&g&!f&e&!a)|(h&!g&f&!e&d&c&b)|(!i&g&!f&!d&!c&b)|(i&!h&g&!e&!b&a)|(i&e&!d&!c&!b&a)|(i&h&!f&e&!d&c)|(!h&g&!d&!c&b&!a)|(!i&g&f&e&!c&b)|(!h&!g&!f&c&b&a)|(i&h&f&d&!c&a)|(!i&g&f&d&c&!a)|(i&h&!e&d&!c&!a)|(!i&f&e&c&!b&a)|(h&f&!e&!d&b&a)|(!h&!g&!f&!d&!c&!b)|(!h&!g&!e&!d&c&a)|(!i&h&!g&f&c&!a)|(!i&h&!g&d&!c&!b)|(!h&!g&!e&d&!c&b)|(h&!g&f&!d&c&!b)|(!f&e&d&c&!b&a)|(i&!h&f&!e&!c&!a)|(i&e&d&c&a)|(i&h&!g&f&a)):((!h&g&!f&!e&d&c&b&a)|(!i&h&!f&e&!d&c&!b&!a)|(!i&!h&!g&!f&!e&c&!b&a)|(i&!h&!g&!f&!e&!d&c&!a)|(i&!h&g&!f&!e&!c&!b&a)|(i&!h&g&f&!e&!d&!c&!a)|(!i&h&g&!f&!e&!c&!b&!a)|(!i&h&g&f&e&d&!c&!a)|(!i&h&!f&e&!d&!c&!b&a)|(!i&!h&!g&f&!e&b&a)|(!i&!h&f&!e&d&b&!a)|(h&f&!e&d&!c&b&!a)|(h&!f&e&d&c&b&a)|(!h&g&!f&!e&c&!b&!a)|(i&h&!f&!e&!c&!b&!a)|(!h&!g&!f&!e&!d&!c&!b)|(!i&h&!g&!d&c&b&a)|(i&g&e&!d&c&b&!a)|(!i&!h&g&!e&!d&c&!a)|(!i&!h&g&e&!d&!c&!a)|(i&f&!e&!d&c&b&a)|(!g&!f&!e&!d&c&b&!a)|(i&h&!g&f&!e&!d&a)|(!i&!h&f&e&d&!c&a)|(i&h&f&e&d&!b&a)|(i&h&!f&!d&c&!b&a)|(!i&!h&!g&f&e&!c&!b)|(i&!h&!g&e&d&c&!b)|(!h&g&f&!e&!d&c&!b)|(h&g&f&!e&d&!c&!b)|(!h&!g&!f&d&!b&!a)|(!i&!h&!f&!c&b&a)|(!i&h&!f&!e&b&!a)|(!i&!h&!g&f&c&!b)|(!i&!f&e&d&!c&!b)|(!h&!g&e&d&c&b)|(!i&g&!f&e&!d&a)|(!i&h&!g&f&e&c)|(!i&h&!e&!c&b&!a)|(i&!h&g&f&!d&!b)|(i&!g&e&!d&!c&!a)|(!i&h&g&!e&!b&a)|(i&h&g&!d&b&a)|(i&h&g&!c&b&!a)|(i&h&g&d&c&!b)|(i&h&g&e&!c&a)|(!i&!h&!g&d&c&b)|(!i&f&d&c&!b)|(g&!f&!d&!c&a));

code[2]<=j?((i&h&!g&!f&!e&!d&!c&!b&a)|(!i&h&!g&!f&!e&d&c&!b&a)|(!i&h&g&f&!e&d&!c&!b&!a)|(!i&h&!g&f&!e&!c&!b&a)|(i&h&!g&!f&e&d&c&b&a)|(!h&!g&!f&!e&!d&!c&b&a)|(!i&h&!g&f&e&!d&!c&b&!a)|(i&!h&!g&f&!e&d&c&b&!a)|(!i&h&!g&f&e&!d&c&!b&!a)|(i&h&g&f&!e&d&c&b&!a)|(i&!h&!g&f&!e&!d&c&b&a)|(!i&h&!g&f&e&d&c&!b&a)|(i&!h&g&e&!d&c&!b&!a)|(i&h&g&f&e&d&!b&!a)|(i&h&!f&!e&d&!c&b&!a)|(i&!g&!f&!e&d&c&b&a)|(h&g&f&e&d&!c&b&!a)|(i&!h&!f&!e&d&!c&!b&a)|(!i&!h&!f&e&d&c&!b&a)|(i&!h&g&f&!e&d&!c&!a)|(!i&h&g&f&!e&c&b&!a)|(!i&h&!g&!f&e&!d&!c&!b)|(i&!h&!g&f&!d&c&!b&a)|(i&!h&!g&f&!d&c&b&!a)|(!i&h&f&!e&!d&!b&a)|(i&!h&!g&f&!e&d&!b&a)|(!i&h&!g&f&d&c&b&!a)|(i&!h&!g&f&!e&!d&!c&!a)|(i&h&g&!f&e&!d&c&!b&a)|(!h&!g&f&e&d&!c&!b&!a)|(!i&!h&!g&f&d&!c&!b&!a)|(!i&h&!g&f&!e&d&c&!a)|(i&g&!f&!e&d&!c&b&a)|(!i&h&g&e&!d&!c&b&a)|(i&!h&g&!f&!d&c&!b&!a)|(i&!h&g&f&!d&c&b&a)|(i&!h&!g&!f&e&!c&!b&a)|(!i&h&g&f&!d&c&!b&a)|(i&!h&g&f&e&d&c&!b)|(i&h&!f&e&!d&!c&b&a)|(i&h&g&f&e&c&b&a)|(!h&!g&!f&!e&!d&c&b&!a)|(!i&h&!g&!f&!e&!d&c&!a)|(h&g&!f&e&d&c&!b&!a)|(i&h&!g&f&!e&!c&b&!a)|(i&!h&!f&!e&!d&c&b&!a)|(i&h&!g&!f&e&d&c&!a)|(!i&!h&g&!e&d&!c&!b&a)|(h&g&f&e&!d&!c&!b&!a)|(i&!g&f&e&d&c&b&a)|(i&h&!g&f&e&d&!c&b)|(h&g&!f&e&!d&b&a)|(!i&!g&f&e&d&!c&!b&!a)|(i&h&!g&f&!e&d&!b&!a)|(!i&!h&!g&f&e&!d&!c&!b)|(i&h&!g&f&!e&d&c&!b)|(!i&h&g&!f&e&!b&!a)|(!i&!h&g&e&!d&b&!a)|(!i&!h&g&!e&c&b&a)|(!h&g&!f&!e&!d&!c&b)|(!i&!h&!g&!f&!d&b&a)|(i&g&f&!e&!d&!c&b)|(!i&!h&g&!e&d&b&!a)|(!h&!f&e&!d&c&!b&!a)|(i&!g&!f&d&c&!b&!a)|(h&!g&!f&e&d&!b&!a)|(!i&h&!g&!f&d&!c&!a)|(!i&h&g&!e&!d&c&!b)|(!i&!h&!g&d&!c&b&a)|(!i&g&f&!e&!d&c&!b)|(i&h&!g&e&!d&c&!b)|(!i&!h&!g&!d&!c&!b&a)|(!i&!h&!g&e&d&!c&b)|(!i&!h&!g&!f&!e&!d&!b)|(!i&h&!g&f&!e&!d&!c)|(i&h&!g&!f&!d&!c&b&!a)|(i&h&g&!f&!d&b&a)|(!i&!h&!g&f&!e&c&!b&a)|(!h&g&e&d&c&b&!a)|(!i&!h&g&!d&!c&b&!a)|(!i&!h&g&!f&!d&!c&!b)|(i&h&e&!d&c&b&!a)|(!i&!h&g&!f&!e&!c&!b)|(!i&h&!g&!f&!e&b&!a)|(!i&!h&f&e&d&!c&!a)|(!h&g&f&e&d&!c&a)|(!i&!h&f&e&!d&!c&a)|(h&!g&!f&!e&!d&b&!a)|(i&h&!g&e&c&!b&!a)|(i&h&f&e&!d&!c&!b)|(!i&h&f&!e&!d&c&a)|(i&!h&f&!e&d&!c&b)):((i&h&!g&!e&d&!c&b&a)|(!i&!h&g&f&d&c&b&!a)|(i&h&!g&!f&e&d&!c&b&a)|(!i&!h&g&!f&!e&d&c&!b&!a)|(i&h&!g&!f&!e&!d&c&!b&!a)|(!i&!h&g&!f&!e&!d&c&b&!a)|(i&!h&g&!f&!e&!d&!c&!b&a)|(i&h&g&!f&!e&d&!c&!b&!a)|(!i&!h&g&f&!e&!d&c&!b&!a)|(!i&h&!g&!f&!e&!d&!c&!b&!a)|(!i&h&g&f&!d&!c&b&a)|(!i&h&g&f&!e&!d&!c&b&!a)|(!i&h&g&f&e&!d&!c&!b&!a)|(i&!h&!f&!e&d&c&!b&a)|(!i&!h&!g&f&e&d&b&!a)|(i&!h&!g&!f&!d&c&b&a)|(i&!h&!g&f&!d&c&b&!a)|(!i&!h&g&f&!e&d&!b&a)|(!i&h&!g&f&d&c&!b&a)|(!i&!h&g&!f&!e&!d&b&a)|(i&!h&g&f&e&d&!c&a)|(!i&!h&!g&f&!d&!c&!b&!a)|(!i&!h&!f&e&d&!c&!b&!a)|(!h&g&!f&e&d&c&!b&a)|(!i&h&!g&!f&e&d&c&b)|(i&!h&!g&!f&e&!d&!c&!a)|(!i&!h&!g&!e&!d&c&!b&a)|(!i&h&g&f&!e&c&!b&!a)|(i&h&g&f&e&!c&b&!a)|(!i&h&!g&f&e&!d&c&!a)|(!i&h&!g&!e&!d&!c&b&a)|(!i&!h&g&f&e&d&!c&!b)|(!i&h&!g&!f&e&!d&!c&!a)|(i&h&g&!e&!d&c&b&a)|(!i&!h&!g&e&!d&c&!b&!a)|(!i&h&g&e&d&c&!b&!a)|(!i&h&!g&f&!e&!d&c&b&a)|(i&h&g&!f&e&!d&!c&!b&!a)|(i&!h&!g&f&!e&d&c&!a)|(!i&!h&!g&!f&d&c&b&!a)|(i&!h&!f&e&d&c&b&a)|(!i&!h&!g&f&!e&d&!c&!a)|(!h&!g&!f&!e&d&!c&!b&!a)|(i&!h&!g&f&e&!d&b&a)|(!i&!g&f&e&d&!c&!b&a)|(i&!h&!g&f&!e&!d&!c&a)|(!i&g&!f&!e&d&!c&!b&a)|(i&!h&!g&!f&!e&!d&!c&b)|(i&h&!g&!e&d&c&b&!a)|(!i&!h&!g&!f&!e&d&!c&a)|(i&!h&g&f&!e&!c&!b&!a)|(i&h&!f&!e&d&!c&b&a)|(h&g&f&e&d&c&b&!a)|(i&!h&!g&e&!d&c&b&!a)|(i&h&!g&!f&e&c&b&!a)|(i&h&!g&f&!e&!d&!b&!a)|(!i&!h&g&f&e&!d&c&b)|(i&!h&g&!f&e&d&!c&!a)|(!i&h&g&!f&e&!d&b&!a)|(!i&h&g&f&!d&!c&!b&a)|(i&!h&g&e&!d&!c&b&a)|(!h&!g&!f&!e&!c&b&a)|(i&!h&!g&f&!c&!b&a)|(i&h&!f&!e&c&b&!a)|(i&g&!f&!e&!d&b&!a)|(i&h&!g&!f&!e&!c&a)|(!h&!g&f&e&d&c&!b)|(!h&!g&!f&e&!d&c&a)|(!i&g&!f&e&!c&b&a)|(!i&g&f&e&d&c&b)|(i&!h&g&f&!d&!b&!a)|(i&h&!f&e&!d&!b&a)|(i&h&!f&e&d&c&!b)|(!i&h&!g&f&e&!d&b)|(!h&!g&f&e&!d&!c&!b)|(i&h&!g&e&c&!b&a)|(i&h&g&!f&!d&c&a)|(!i&h&g&!f&d&!c&b)|(h&!g&e&d&!c&!b&!a)|(!i&h&g&!e&d&!c&a)|(!i&h&g&f&e&d&c)|(i&!h&g&e&c&!b&!a)|(h&g&!e&!d&!c&!b&a)|(!i&h&g&!e&!d&!c&!b)|(h&!g&!f&e&d&c&!b&a)|(i&g&f&e&d&!c&b)|(!i&g&f&!e&!d&!c&a)|(!i&h&!g&!f&!e&c&!a)|(i&h&g&!f&e&b&a)|(i&!h&!g&!d&!c&!b&a)|(h&g&!f&e&!d&c&!b));

code[1]<=j?((!i&h&g&f&e&d&!c&!b&a)|(i&h&!g&!f&e&d&c&b&a)|(!h&!g&!f&!e&!d&!c&b&a)|(!i&h&!g&f&e&!d&!c&b&!a)|(i&!h&!g&f&!e&d&c&b&!a)|(i&h&!g&f&e&!d&c&!b&a)|(!i&h&!g&f&e&!d&c&!b&!a)|(!i&g&!f&e&!d&!c&!b&!a)|(i&!h&g&!f&!e&d&!c&!a)|(i&!h&!f&e&d&c&!b&a)|(i&h&!g&!f&d&!c&!b&a)|(!i&g&f&!e&!d&c&b&a)|(i&h&!g&!f&e&!c&!b&!a)|(!i&!g&!f&e&d&c&!b&a)|(i&h&f&!e&d&c&b&a)|(!i&h&!g&!f&e&!d&c&b)|(h&!f&!e&!d&c&!b&a)|(!i&h&!g&f&e&c&b&a)|(!i&!h&!g&!e&!d&!c&b&a)|(i&h&!g&f&!d&!c&!b&!a)|(!i&h&f&!e&d&c&b&!a)|(i&!g&f&!e&d&c&!b&!a)|(i&h&g&!f&e&!d&c&!b&a)|(i&g&!f&!e&d&!c&b&a)|(!i&h&g&e&!d&!c&b&a)|(i&!h&g&!f&!d&c&!b&!a)|(i&!h&g&f&!d&c&b&a)|(i&!h&g&e&d&!c&b&a)|(i&!h&!g&!f&e&!c&!b&a)|(!i&h&g&f&!d&c&!b&a)|(i&g&f&e&!d&!c&!b&a)|(i&!h&g&f&e&d&c&!b)|(!h&!g&!f&!e&!d&c&b&!a)|(!i&h&!g&!f&!e&!d&c&!a)|(i&h&!g&f&!e&!c&b&!a)|(i&!h&!g&e&!d&!c&b&!a)|(!i&h&g&f&!e&!d&!b&!a)|(i&!h&g&f&!e&d&c&!b)|(h&!g&f&e&d&c&!b&!a)|(h&!g&f&!e&d&!c&!b&a)|(i&h&g&!f&!d&c&b)|(i&h&g&e&!d&b&!a)|(!h&!g&f&!e&d&c&!b&!a)|(h&g&!f&!e&c&!b&a)|(i&g&!f&!e&!d&!c&!b)|(h&g&e&!d&c&b&!a)|(i&!h&g&!e&d&b&!a)|(!h&g&f&e&!d&c&a)|(!i&!g&!f&d&!c&b&a)|(i&h&g&f&e&d&c)|(h&g&!e&d&!c&b&!a)|(i&!h&!g&!f&!d&b&!a)|(i&!h&f&e&d&!c&a)|(i&!h&f&e&!d&c&a)|(!i&!h&g&!f&!e&!d&!b)|(i&g&f&!e&!d&!b&!a)|(h&!g&!f&!e&!c&b&a)|(!i&!h&g&f&!e&b&!a)|(!i&!h&!g&!f&c&!b&a)|(!i&!h&!f&e&d&!c&!b)|(!g&f&e&d&!c&b&a)|(!i&!h&!e&d&c&b&a)|(!i&f&!e&!d&!c&!b&a)|(i&!h&!g&!d&c&!b&!a)|(!i&!h&f&!e&d&c&a)|(!h&!g&f&e&d&b&!a)|(i&h&!g&f&!e&!d&b)|(!i&!h&!g&f&e&c&!a)|(!i&!g&f&e&!d&!c&!b)|(i&h&!g&!f&!d&!c&b&!a)|(i&h&g&!f&!d&b&a)|(!i&!h&!g&f&!e&c&!b&a)|(!h&g&e&d&c&b&!a)|(!i&!h&g&!d&!c&b&!a)|(!i&!h&g&!f&!d&!c&!b)|(i&h&e&!d&c&b&!a)|(!i&!h&g&!f&!e&!c&!b)|(!i&h&!g&!f&!e&b&!a)|(!i&!h&f&e&d&!c&!a)|(!i&!h&g&f&e&!c&b)|(g&f&!e&!c&b&!a)|(!h&!g&!f&e&c&!b)|(!i&!e&d&!c&!b&!a)):((i&!h&g&!f&e&!c&!b&!a)|(i&h&!g&!f&e&d&!c&b&a)|(!i&!h&g&!f&!e&d&c&!b&!a)|(!i&h&!g&!f&!e&d&c&b&a)|(i&h&!g&!f&!e&!d&c&!b&!a)|(!i&!h&g&!f&!e&!d&c&b&!a)|(i&!h&g&!f&!e&!d&!c&!b&a)|(i&!h&g&f&e&d&c&b&a)|(i&h&g&!f&!e&d&!c&!b&!a)|(!i&!h&g&f&!e&!d&c&!b&!a)|(!i&h&!g&!f&!e&!d&!c&!b&!a)|(!i&h&g&f&!d&!c&b&a)|(!i&h&g&f&e&!d&!c&!b&!a)|(!h&!g&f&!e&d&c&b&a)|(i&f&e&d&!c&b&!a)|(i&!h&f&!e&!d&!c&b&a)|(!h&!g&f&!e&!d&!c&b&!a)|(i&!h&!g&!f&!d&c&b&!a)|(!i&h&f&!e&d&!c&b&a)|(!i&!h&!g&!f&!d&c&b&a)|(i&h&!g&f&d&!c&!b&!a)|(!i&h&!f&!e&d&c&!b&!a)|(i&!h&g&!e&d&c&b&!a)|(i&g&f&!e&!d&!c&!b&!a)|(!i&h&!g&f&e&d&!c&b)|(!i&h&f&!e&!d&!c&!b&a)|(i&!h&g&!e&!d&c&b&a)|(i&!h&!g&!f&e&!d&c&!b)|(!i&!h&g&f&e&!c&!b&a)|(!h&g&f&e&!d&!c&!b&a)|(i&h&!g&f&e&!d&c&!b)|(i&!h&g&!f&e&!d&!c&!a)|(!i&h&g&e&!d&!c&b&!a)|(!i&h&!g&f&!e&!d&c&b&a)|(i&h&g&!f&e&!d&!c&!b&!a)|(i&!h&!g&f&!e&d&c&!a)|(!i&!h&!g&!f&d&c&b&!a)|(i&!h&!f&e&d&c&b&a)|(!i&!h&!g&f&!e&d&!c&!a)|(!h&!g&!f&!e&d&!c&!b&!a)|(i&!h&!g&f&e&!d&b&a)|(!i&!g&f&e&d&!c&!b&a)|(i&!h&!g&f&!e&!d&!c&a)|(!i&g&!f&!e&d&!c&!b&a)|(i&!h&!g&!f&!e&!d&!c&b)|(i&h&!g&!e&d&c&b&!a)|(!h&!g&f&!e&d&c&!b&!a)|(i&!h&g&f&!e&!c&!b&!a)|(i&!h&!f&e&d&!c&b&a)|(h&g&f&e&d&c&b&!a)|(i&!h&!g&e&!d&c&b&!a)|(!i&g&!f&!e&!d&!c&b&a)|(!i&!h&g&f&e&!d&c&b)|(!i&h&g&f&!e&d&!b&!a)|(i&h&g&!f&!e&d&!c&b)|(i&h&!f&e&!d&c&b&!a)|(!i&!h&!g&!f&e&!d&!c&!a)|(!i&!h&f&e&!d&!c&!b&!a)|(h&g&!f&!e&!d&c&!b&a)|(!i&h&g&!f&e&d&!c&!b)|(i&!g&f&!e&d&b&a)|(!h&!f&!e&d&!c&b&!a)|(!i&!g&!f&!e&d&!c&!a)|(!i&!h&!f&d&!c&b&!a)|(i&g&f&d&c&!b&a)|(!i&h&f&!e&c&b&!a)|(!i&!h&!g&!f&e&!b&a)|(i&!h&!g&!e&c&!b&a)|(!h&g&f&!d&c&b&a)|(!i&h&!g&!f&!e&d&!b)|(i&h&f&!d&c&!b&a)|(!h&!g&e&d&!c&!b&a)|(!h&g&!e&d&c&!b&a)|(i&h&g&!f&d&c&b)|(!i&!g&e&!d&c&b&!a)|(i&h&!g&!f&e&!d&b)|(!i&!h&!f&!e&!d&!c&!b)|(h&g&f&!e&!d&c&b)|(h&g&!e&d&!c&!b&a)|(!i&!h&g&e&!d&b&a)|(!i&!h&g&e&c&!b&!a)|(h&g&e&!d&c&!b&a)|(h&!g&!f&e&d&c&!b&a)|(i&g&f&e&d&!c&b)|(!i&g&f&!e&!d&!c&a)|(!h&!g&!f&e&d&c&!a)|(i&!g&e&!d&!c&b&a)|(i&h&!g&e&d&!c&!a)|(h&g&!f&e&!d&c&!b)|(g&!f&e&d&c&!a)|(i&h&g&f&e&d));

code[0]<=j?((!i&!h&!g&f&!e&!d&c&b&!a)|(i&h&!g&f&e&!d&c&!b&a)|(i&h&g&f&!e&d&c&b&!a)|(i&!h&!g&f&!e&!d&c&b&a)|(!i&h&!g&f&e&d&c&!b&a)|(!i&g&!f&e&!d&c&b&!a)|(i&!h&!f&e&d&c&b&!a)|(h&g&!f&!e&!d&c&!b&!a)|(i&h&g&f&!e&!c&!b&a)|(!i&!h&g&e&d&!c&!b&!a)|(!h&g&!f&!e&d&c&!b&!a)|(!i&!h&g&!e&!d&c&!b&a)|(i&h&g&f&!e&!d&c&b)|(i&h&g&!f&e&!d&c&!b&a)|(!i&!h&g&f&!e&d&c&b)|(!i&!g&!f&!e&d&!c&!b&!a)|(!i&!h&!g&!f&e&d&c)|(i&h&g&!f&e&d&b&a)|(!i&!h&!g&f&e&d&b&!a)|(!i&!h&!g&!e&!d&c&!b&!a)|(!g&f&!e&d&!c&b&!a)|(!h&!g&!f&e&d&!c&b&a)|(!i&!h&!g&!f&e&!d&b&!a)|(!i&h&!g&e&d&!c&b&!a)|(!h&!g&f&!e&!d&!c&!b&a)|(i&!h&g&e&d&!c&b&a)|(i&g&f&e&!d&!c&!b&a)|(i&h&!f&e&!d&!c&b&a)|(i&h&g&f&e&c&b&a)|(h&g&!f&e&d&c&!b&!a)|(i&!h&!g&e&!d&!c&b&!a)|(i&!h&!f&!e&!d&c&b&!a)|(i&h&!g&!f&e&d&c&!a)|(!i&h&g&f&!e&!d&!b&!a)|(!i&!h&g&!e&d&!c&!b&a)|(i&!h&g&f&!e&d&c&!b)|(h&g&f&e&!d&!c&!b&!a)|(i&!g&f&e&d&c&b&a)|(i&h&!g&f&e&d&!c&b)|(h&!g&f&e&d&c&!b&!a)|(h&!g&f&!e&d&!c&!b&a)|(!i&!g&f&e&d&!c&!b&!a)|(i&h&!g&f&!e&d&!b&!a)|(!h&!g&f&!e&d&c&!b&!a)|(!i&!h&!g&f&e&!d&!c&!b)|(i&h&!g&f&!e&d&c&!b)|(!h&g&!f&e&!d&b&a)|(i&h&g&!f&e&!c&!b)|(!i&h&g&!f&!e&!c&a)|(!i&g&!e&!d&!c&b&a)|(i&g&f&d&!c&b&!a)|(i&!h&g&!f&!e&d&c)|(i&!h&g&!f&!e&!c&!b)|(!i&h&g&!f&!e&c&b)|(!h&g&f&!d&!c&b&a)|(i&!h&f&e&d&b&a)|(i&!f&!e&!d&!c&!b&!a)|(!i&!g&!f&e&c&!b&a)|(i&!h&!f&e&!d&c&!b)|(i&!g&!f&!e&c&!b&a)|(!h&!f&e&!d&!c&!b&!a)|(i&!h&g&f&d&!b&!a)|(i&!h&!g&!f&e&!d&!c)|(!i&!h&g&!e&!d&!c&!a)|(!i&h&!g&!f&!e&!d&a)|(i&h&f&e&!d&!b&!a)|(i&!g&e&d&!c&!b&!a)|(i&!h&!f&!e&d&c&!b)|(!i&!h&!g&!f&d&c&b)|(h&!g&f&e&!d&b&!a)|(h&f&!e&d&!c&b&!a)|(!i&h&!g&!e&!c&b&!a)|(!i&!h&f&e&!d&c&!b)|(!i&h&f&!e&c&!b&!a)|(!i&h&!g&!e&d&!b&!a)|(i&h&!g&!f&!d&!c&b&!a)|(h&g&f&d&c&!b&a)|(h&!g&e&!d&!c&b&a)|(i&h&!g&!e&!d&b&a)|(!i&h&g&f&e&d&c)|(i&!h&!g&!e&d&b&a)|(!i&h&!g&!f&!e&!c&!a)|(!i&!h&!g&f&!e&c&!b&a)|(h&!g&f&!e&d&c&b)|(!i&!h&g&f&e&!c&b)|(!h&g&f&e&d&!c&a)|(!i&!h&f&e&!d&!c&a)|(h&!g&!f&!e&!d&b&!a)|(i&h&!g&e&c&!b&!a)|(i&h&f&e&!d&!c&!b)|(!i&h&f&!e&!d&c&a)|(i&!h&f&!e&d&!c&b)|(i&g&!f&d&c&!b)|(!i&h&!f&e&d&a)|(!i&h&g&f&e&a)|(i&h&!f&e&d&!c)|(i&!g&!f&!e&!c&b)|(h&!f&!e&!d&!c&b)|(!i&!h&!g&e&c&a)|(!i&g&f&d&!c&!b)|(!i&!h&f&e&!b&a)|(!f&e&d&c&!b&a)|(i&!h&f&!e&!c&!a)):((!i&h&!g&!f&!e&d&c&b&a)|(i&!h&g&f&e&d&c&b&a)|(!i&h&g&f&!e&!d&!c&b&!a)|(i&g&f&!e&d&!c&b&a)|(!i&!h&g&!f&e&d&b&a)|(i&!h&g&!f&!d&c&b&!a)|(!i&h&!g&f&!d&c&!b&!a)|(i&!h&g&!e&d&c&!b&!a)|(i&!h&g&e&d&c&b&!a)|(h&!g&!f&e&!d&!c&!b&!a)|(i&h&g&f&!d&c&!b&!a)|(!i&h&!g&e&d&c&!b&!a)|(!i&!h&g&e&d&c&!b&!a)|(i&h&g&f&e&!d&c&!a)|(i&!h&g&!e&!d&!c&!b&!a)|(!i&h&!g&e&!d&c&!b&a)|(!i&!h&g&!f&e&!d&!c&!b)|(!i&h&!g&f&!e&!d&c&b&a)|(!i&!h&!g&!f&!e&c&!b&a)|(i&!h&!g&!f&!e&!d&c&!a)|(i&!h&g&!f&!e&!c&!b&a)|(i&h&g&!f&e&!d&!c&!b&!a)|(i&!h&g&f&!e&!d&!c&!a)|(!i&h&g&!f&!e&!c&!b&!a)|(!i&h&g&f&e&d&!c&!a)|(!i&h&!f&e&!d&!c&!b&a)|(!h&!g&f&!e&d&c&!b&!a)|(!i&!h&!g&!f&!e&d&!c&a)|(i&h&!f&!e&d&!c&b&a)|(i&!h&!f&e&d&!c&b&a)|(i&h&!g&!f&e&c&b&!a)|(i&h&!g&f&!e&!d&!b&!a)|(!i&g&!f&!e&!d&!c&b&a)|(!i&h&g&f&!e&d&!b&!a)|(i&!h&g&!f&e&d&!c&!a)|(i&h&g&!f&!e&d&!c&b)|(i&h&!f&e&!d&c&b&!a)|(!i&!h&!g&!f&e&!d&!c&!a)|(!i&!h&f&e&!d&!c&!b&!a)|(h&g&!f&!e&!d&c&!b&a)|(!i&h&g&!f&e&!d&b&!a)|(!i&h&g&f&!d&!c&!b&a)|(i&!h&g&e&!d&!c&b&a)|(!i&h&g&!f&e&d&!c&!b)|(i&!h&!g&f&!e&d&!a)|(i&f&!e&d&c&!b&a)|(!i&!h&!g&f&!e&c&b)|(i&!g&f&e&d&!c&b)|(!i&g&f&!e&d&c&b)|(!i&!h&!g&!f&!e&!d&!a)|(i&h&g&f&!e&b&a)|(i&h&!g&f&!e&d&c)|(!i&!h&f&!e&!c&!b&!a)|(i&!h&g&f&d&c&!a)|(i&h&!g&!f&d&!c&!a)|(i&h&!g&f&!c&!b&a)|(i&g&!f&!e&!d&!b&a)|(!i&h&!g&!f&d&!c&b)|(!i&!g&f&e&!d&!c&!a)|(!i&!h&!g&d&!c&!b&a)|(g&!f&e&!d&c&b&a)|(!i&f&e&!d&c&!b&!a)|(h&!g&e&d&c&b&a)|(i&!h&g&!f&e&!c&a)|(h&g&f&e&!c&b&a)|(i&h&!g&!e&!d&c&a)|(!i&h&!g&!e&d&!c&b)|(!i&h&!f&!e&!d&!c&b)|(!i&h&g&!e&c&b&a)|(h&!g&f&e&!d&!c&b)|(i&h&!g&!d&!c&b&!a)|(!i&!h&g&!e&!d&!b&a)|(i&h&!f&e&!d&!c&b)|(i&g&f&e&!d&!c&!b)|(i&h&g&e&d&!b&!a)|(h&g&e&d&c&!b&a)|(!i&h&g&e&!d&b&a)|(h&!g&!f&e&d&c&!b&a)|(i&f&!e&!d&c&b&a)|(!g&!f&!e&!d&c&b&!a)|(i&h&!g&f&!e&!d&a)|(!i&!h&f&e&d&!c&a)|(i&h&f&e&d&!b&a)|(i&h&!f&!d&c&!b&a)|(!i&!h&!g&f&e&!c&!b)|(i&!h&!g&e&d&c&!b)|(!h&g&f&!e&!d&c&!b)|(h&g&f&!e&d&!c&!b)|(!h&!g&!f&e&d&c&!a)|(!i&h&!g&!f&!e&c&!a)|(i&h&g&!f&e&b&a)|(i&!g&e&!d&!c&b&a)|(i&!h&!g&!d&!c&!b&a)|(i&h&!g&e&d&!c&!a)|(!i&!g&f&!e&d&a)|(!h&!g&!f&d&b&!a)|(i&h&!g&f&e&b)|(i&h&!f&d&c&!b)|(!i&!h&!g&d&c&b));
		end

	end

	decoder decoder(.code(code), .segments(io_out));

endmodule
